VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3520.000 BY 3710.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1504.200 3520.000 1504.800 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2688.790 3706.000 2689.070 3710.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2297.330 3706.000 2297.610 3710.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 3706.000 1906.610 3710.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 3706.000 1515.610 3710.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 3706.000 1124.610 3710.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 3706.000 733.150 3710.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 3706.000 342.150 3710.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3674.760 4.000 3675.360 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3400.040 4.000 3400.640 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3125.320 4.000 3125.920 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1784.360 3520.000 1784.960 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2850.600 4.000 2851.200 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2575.880 4.000 2576.480 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2301.160 4.000 2301.760 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2026.440 4.000 2027.040 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1476.320 4.000 1476.920 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1201.600 4.000 1202.200 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.880 4.000 927.480 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2064.520 3520.000 2065.120 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2344.680 3520.000 2345.280 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2624.160 3520.000 2624.760 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2904.320 3520.000 2904.920 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3184.480 3520.000 3185.080 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3464.640 3520.000 3465.240 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3470.790 3706.000 3471.070 3710.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3079.790 3706.000 3080.070 3710.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 34.720 3520.000 35.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2414.720 3520.000 2415.320 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2694.200 3520.000 2694.800 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2974.360 3520.000 2974.960 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3254.520 3520.000 3255.120 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3534.680 3520.000 3535.280 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3372.810 3706.000 3373.090 3710.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.810 3706.000 2982.090 3710.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2590.810 3706.000 2591.090 3710.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.810 3706.000 2200.090 3710.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.810 3706.000 1809.090 3710.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 244.160 3520.000 244.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 3706.000 1417.630 3710.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 3706.000 1026.630 3710.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 3706.000 635.630 3710.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 3706.000 244.630 3710.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3606.080 4.000 3606.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3331.360 4.000 3331.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3056.640 4.000 3057.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2781.920 4.000 2782.520 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2507.200 4.000 2507.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2232.480 4.000 2233.080 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 454.280 3520.000 454.880 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1957.760 4.000 1958.360 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1682.360 4.000 1682.960 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.920 4.000 1133.520 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 664.400 3520.000 665.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 874.520 3520.000 875.120 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1084.640 3520.000 1085.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1294.080 3520.000 1294.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1574.240 3520.000 1574.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1854.400 3520.000 1855.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2134.560 3520.000 2135.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 174.120 3520.000 174.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2554.120 3520.000 2554.720 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2834.280 3520.000 2834.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3114.440 3520.000 3115.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3394.600 3520.000 3395.200 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3674.760 3520.000 3675.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3177.310 3706.000 3177.590 3710.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.310 3706.000 2786.590 3710.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.310 3706.000 2395.590 3710.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.310 3706.000 2004.590 3710.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.850 3706.000 1613.130 3710.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 384.240 3520.000 384.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 3706.000 1222.130 3710.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 3706.000 831.130 3710.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 3706.000 440.130 3710.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 3706.000 49.130 3710.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3468.720 4.000 3469.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3194.000 4.000 3194.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2919.280 4.000 2919.880 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2644.560 4.000 2645.160 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2369.840 4.000 2370.440 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2095.120 4.000 2095.720 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 594.360 3520.000 594.960 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.720 4.000 1820.320 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1545.000 4.000 1545.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 995.560 4.000 996.160 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 804.480 3520.000 805.080 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1014.600 3520.000 1015.200 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1224.720 3520.000 1225.320 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1434.160 3520.000 1434.760 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1714.320 3520.000 1714.920 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1994.480 3520.000 1995.080 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2274.640 3520.000 2275.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 104.080 3520.000 104.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2484.760 3520.000 2485.360 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2764.240 3520.000 2764.840 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3044.400 3520.000 3045.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3324.560 3520.000 3325.160 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 3604.720 3520.000 3605.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3275.290 3706.000 3275.570 3710.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2884.290 3706.000 2884.570 3710.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.830 3706.000 2493.110 3710.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.830 3706.000 2102.110 3710.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.830 3706.000 1711.110 3710.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 314.200 3520.000 314.800 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 3706.000 1320.110 3710.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 3706.000 929.110 3710.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 3706.000 537.650 3710.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 3706.000 146.650 3710.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3537.400 4.000 3538.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3262.680 4.000 3263.280 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2987.960 4.000 2988.560 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2713.240 4.000 2713.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2438.520 4.000 2439.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2163.800 4.000 2164.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 524.320 3520.000 524.920 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1889.080 4.000 1889.680 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.680 4.000 1614.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1338.960 4.000 1339.560 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 734.440 3520.000 735.040 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 944.560 3520.000 945.160 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1154.680 3520.000 1155.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1364.120 3520.000 1364.720 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1644.280 3520.000 1644.880 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 1924.440 3520.000 1925.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3516.000 2204.600 3520.000 2205.200 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2895.790 0.000 2896.070 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2917.410 0.000 2917.690 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2938.570 0.000 2938.850 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2960.190 0.000 2960.470 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.350 0.000 2981.630 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3002.970 0.000 3003.250 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3024.130 0.000 3024.410 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3045.750 0.000 3046.030 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3066.910 0.000 3067.190 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3088.530 0.000 3088.810 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3109.690 0.000 3109.970 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3131.310 0.000 3131.590 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3152.470 0.000 3152.750 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3173.630 0.000 3173.910 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3195.250 0.000 3195.530 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3216.410 0.000 3216.690 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3238.030 0.000 3238.310 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3259.190 0.000 3259.470 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3280.810 0.000 3281.090 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3301.970 0.000 3302.250 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 0.000 993.970 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3323.590 0.000 3323.870 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3344.750 0.000 3345.030 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3366.370 0.000 3366.650 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3387.530 0.000 3387.810 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3409.150 0.000 3409.430 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3430.310 0.000 3430.590 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3451.930 0.000 3452.210 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3473.090 0.000 3473.370 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 0.000 1015.130 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 0.000 1036.750 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 0.000 1057.910 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.410 0.000 1100.690 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.130 0.000 1207.410 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 0.000 1229.030 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 0.000 1250.190 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.690 0.000 1292.970 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.090 0.000 1357.370 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.190 0.000 1442.470 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.810 0.000 1464.090 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 0.000 1485.250 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 0.000 1506.870 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.370 0.000 1549.650 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 0.000 1570.810 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.150 0.000 1592.430 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 0.000 1635.210 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 0.000 1656.370 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 0.000 1699.150 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.490 0.000 1720.770 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.270 0.000 1763.550 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 0.000 1784.710 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.590 0.000 1805.870 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.210 0.000 1827.490 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 0.000 1848.650 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.990 0.000 1870.270 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.150 0.000 1891.430 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 0.000 1913.050 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.930 0.000 1934.210 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.550 0.000 1955.830 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.710 0.000 1976.990 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.330 0.000 1998.610 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.490 0.000 2019.770 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 0.000 2041.390 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.270 0.000 2062.550 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.890 0.000 2084.170 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.050 0.000 2105.330 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.210 0.000 2126.490 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.610 0.000 2190.890 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2211.770 0.000 2212.050 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2233.390 0.000 2233.670 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.550 0.000 2254.830 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.170 0.000 2276.450 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2297.330 0.000 2297.610 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.950 0.000 2319.230 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.110 0.000 2340.390 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.730 0.000 2362.010 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 0.000 2383.170 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.510 0.000 2404.790 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.670 0.000 2425.950 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.290 0.000 2447.570 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2468.450 0.000 2468.730 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.610 0.000 2489.890 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.230 0.000 2511.510 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.390 0.000 2532.670 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.010 0.000 2554.290 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.170 0.000 2575.450 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.790 0.000 2597.070 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2617.950 0.000 2618.230 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2639.570 0.000 2639.850 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.730 0.000 2661.010 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.350 0.000 2682.630 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.510 0.000 2703.790 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2725.130 0.000 2725.410 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2746.290 0.000 2746.570 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.910 0.000 2768.190 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2789.070 0.000 2789.350 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.690 0.000 2810.970 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2831.850 0.000 2832.130 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2853.010 0.000 2853.290 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.630 0.000 2874.910 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 0.000 765.810 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2903.150 0.000 2903.430 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2924.310 0.000 2924.590 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2945.930 0.000 2946.210 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2967.090 0.000 2967.370 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2988.710 0.000 2988.990 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3009.870 0.000 3010.150 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3031.490 0.000 3031.770 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3052.650 0.000 3052.930 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3074.270 0.000 3074.550 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3095.430 0.000 3095.710 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3117.050 0.000 3117.330 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3138.210 0.000 3138.490 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3159.830 0.000 3160.110 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3180.990 0.000 3181.270 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3202.150 0.000 3202.430 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3223.770 0.000 3224.050 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3244.930 0.000 3245.210 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3266.550 0.000 3266.830 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3287.710 0.000 3287.990 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3309.330 0.000 3309.610 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3330.490 0.000 3330.770 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3352.110 0.000 3352.390 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3373.270 0.000 3373.550 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3394.890 0.000 3395.170 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3416.050 0.000 3416.330 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3437.670 0.000 3437.950 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3458.830 0.000 3459.110 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3480.450 0.000 3480.730 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.310 0.000 1107.590 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 0.000 1171.990 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.870 0.000 1193.150 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 0.000 1214.770 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 0.000 1300.330 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.210 0.000 1321.490 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 0.000 1385.890 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.770 0.000 1407.050 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 0.000 1449.830 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.710 0.000 1470.990 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 0.000 1535.390 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.270 0.000 1556.550 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 0.000 1599.330 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.670 0.000 1620.950 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.830 0.000 1642.110 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.450 0.000 1663.730 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 0.000 1684.890 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 0.000 1706.510 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.390 0.000 1727.670 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.010 0.000 1749.290 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.170 0.000 1770.450 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.110 0.000 1834.390 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.730 0.000 1856.010 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.890 0.000 1877.170 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.510 0.000 1898.790 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 0.000 1919.950 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.290 0.000 1941.570 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.450 0.000 1962.730 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.070 0.000 1984.350 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.230 0.000 2005.510 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.850 0.000 2027.130 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 0.000 2048.290 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.790 0.000 2091.070 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 0.000 2112.690 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.570 0.000 2133.850 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.730 0.000 2155.010 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.350 0.000 2176.630 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.510 0.000 2197.790 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.130 0.000 2219.410 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.290 0.000 2240.570 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2261.910 0.000 2262.190 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.690 0.000 2304.970 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.850 0.000 2326.130 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.470 0.000 2347.750 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.630 0.000 2368.910 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.250 0.000 2390.530 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.410 0.000 2411.690 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.030 0.000 2433.310 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.190 0.000 2454.470 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.350 0.000 2475.630 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.970 0.000 2497.250 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 0.000 2518.410 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2539.750 0.000 2540.030 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.910 0.000 2561.190 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.530 0.000 2582.810 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.690 0.000 2603.970 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.310 0.000 2625.590 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.470 0.000 2646.750 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.090 0.000 2668.370 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2689.250 0.000 2689.530 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2710.870 0.000 2711.150 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.030 0.000 2732.310 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.650 0.000 2753.930 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.810 0.000 2775.090 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2796.430 0.000 2796.710 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2817.590 0.000 2817.870 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2838.750 0.000 2839.030 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2860.370 0.000 2860.650 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.530 0.000 2881.810 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 0.000 958.090 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.050 0.000 2910.330 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2931.670 0.000 2931.950 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2952.830 0.000 2953.110 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2974.450 0.000 2974.730 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2995.610 0.000 2995.890 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3017.230 0.000 3017.510 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3038.390 0.000 3038.670 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3060.010 0.000 3060.290 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3081.170 0.000 3081.450 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3102.790 0.000 3103.070 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 0.000 986.610 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3123.950 0.000 3124.230 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3145.570 0.000 3145.850 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3166.730 0.000 3167.010 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3187.890 0.000 3188.170 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3209.510 0.000 3209.790 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3230.670 0.000 3230.950 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3252.290 0.000 3252.570 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3273.450 0.000 3273.730 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3295.070 0.000 3295.350 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3316.230 0.000 3316.510 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3337.850 0.000 3338.130 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3359.010 0.000 3359.290 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3380.630 0.000 3380.910 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3401.790 0.000 3402.070 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3423.410 0.000 3423.690 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3444.570 0.000 3444.850 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3466.190 0.000 3466.470 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3487.350 0.000 3487.630 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 0.000 1114.950 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.790 0.000 1286.070 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 0.000 1307.230 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 0.000 1328.850 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 0.000 1371.630 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 0.000 1392.790 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.450 0.000 1456.730 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.230 0.000 1499.510 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.850 0.000 1521.130 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.010 0.000 1542.290 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 0.000 1585.070 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 0.000 1606.690 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.190 0.000 1649.470 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.350 0.000 1670.630 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 0.000 1735.030 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.910 0.000 1756.190 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.070 0.000 1777.350 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.690 0.000 1798.970 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 0.000 1820.130 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.470 0.000 1841.750 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.630 0.000 1862.910 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.250 0.000 1884.530 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.030 0.000 1927.310 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.810 0.000 1970.090 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.970 0.000 1991.250 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 0.000 2012.870 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.750 0.000 2034.030 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.370 0.000 2055.650 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.530 0.000 2076.810 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.150 0.000 2098.430 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.310 0.000 2119.590 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.470 0.000 2140.750 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.090 0.000 2162.370 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 0.000 2183.530 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.870 0.000 2205.150 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.030 0.000 2226.310 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 0.000 901.050 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.810 0.000 2269.090 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.430 0.000 2290.710 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.590 0.000 2311.870 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.210 0.000 2333.490 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2354.370 0.000 2354.650 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.990 0.000 2376.270 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2397.150 0.000 2397.430 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2418.770 0.000 2419.050 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.930 0.000 2440.210 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.550 0.000 2461.830 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 0.000 922.670 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.710 0.000 2482.990 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2503.870 0.000 2504.150 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2525.490 0.000 2525.770 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2546.650 0.000 2546.930 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2568.270 0.000 2568.550 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.430 0.000 2589.710 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.050 0.000 2611.330 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.210 0.000 2632.490 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2653.830 0.000 2654.110 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.990 0.000 2675.270 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.610 0.000 2696.890 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.770 0.000 2718.050 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.390 0.000 2739.670 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2760.550 0.000 2760.830 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2782.170 0.000 2782.450 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.330 0.000 2803.610 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2824.490 0.000 2824.770 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2846.110 0.000 2846.390 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2867.270 0.000 2867.550 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2888.890 0.000 2889.170 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3494.710 0.000 3494.990 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3501.610 0.000 3501.890 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3508.970 0.000 3509.250 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3515.870 0.000 3516.150 4.000 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3424.020 -9.320 3427.020 3716.680 ;
    END
  END vccd1
  PIN vccd1.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3244.020 -9.320 3247.020 3716.680 ;
    END
  END vccd1.extra1
  PIN vccd1.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3064.020 3669.800 3067.020 3716.680 ;
    END
  END vccd1.extra2
  PIN vccd1.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2884.020 3669.800 2887.020 3716.680 ;
    END
  END vccd1.extra3
  PIN vccd1.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2704.020 3669.800 2707.020 3716.680 ;
    END
  END vccd1.extra4
  PIN vccd1.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2524.020 3669.800 2527.020 3716.680 ;
    END
  END vccd1.extra5
  PIN vccd1.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2344.020 3669.800 2347.020 3716.680 ;
    END
  END vccd1.extra6
  PIN vccd1.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2164.020 3669.800 2167.020 3716.680 ;
    END
  END vccd1.extra7
  PIN vccd1.extra8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1984.020 3669.800 1987.020 3716.680 ;
    END
  END vccd1.extra8
  PIN vccd1.extra9
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1804.020 3669.800 1807.020 3716.680 ;
    END
  END vccd1.extra9
  PIN vccd1.extra10
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1624.020 3669.800 1627.020 3716.680 ;
    END
  END vccd1.extra10
  PIN vccd1.extra11
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1444.020 3669.800 1447.020 3716.680 ;
    END
  END vccd1.extra11
  PIN vccd1.extra12
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1264.020 3669.800 1267.020 3716.680 ;
    END
  END vccd1.extra12
  PIN vccd1.extra13
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1084.020 3669.800 1087.020 3716.680 ;
    END
  END vccd1.extra13
  PIN vccd1.extra14
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 904.020 3669.800 907.020 3716.680 ;
    END
  END vccd1.extra14
  PIN vccd1.extra15
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 724.020 3669.800 727.020 3716.680 ;
    END
  END vccd1.extra15
  PIN vccd1.extra16
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 544.020 3669.800 547.020 3716.680 ;
    END
  END vccd1.extra16
  PIN vccd1.extra17
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 364.020 3669.800 367.020 3716.680 ;
    END
  END vccd1.extra17
  PIN vccd1.extra18
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.020 -9.320 187.020 3716.680 ;
    END
  END vccd1.extra18
  PIN vccd1.extra19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.020 -9.320 7.020 3716.680 ;
    END
  END vccd1.extra19
  PIN vccd1.extra20
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3526.900 -4.620 3529.900 3711.980 ;
    END
  END vccd1.extra20
  PIN vccd1.extra21
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3711.980 ;
    END
  END vccd1.extra21
  PIN vccd1.extra22
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3064.020 -9.320 3067.020 430.000 ;
    END
  END vccd1.extra22
  PIN vccd1.extra23
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2884.020 -9.320 2887.020 430.000 ;
    END
  END vccd1.extra23
  PIN vccd1.extra24
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2704.020 -9.320 2707.020 430.000 ;
    END
  END vccd1.extra24
  PIN vccd1.extra25
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2524.020 -9.320 2527.020 430.000 ;
    END
  END vccd1.extra25
  PIN vccd1.extra26
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2344.020 -9.320 2347.020 430.000 ;
    END
  END vccd1.extra26
  PIN vccd1.extra27
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2164.020 -9.320 2167.020 430.000 ;
    END
  END vccd1.extra27
  PIN vccd1.extra28
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1984.020 -9.320 1987.020 430.000 ;
    END
  END vccd1.extra28
  PIN vccd1.extra29
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1804.020 -9.320 1807.020 430.000 ;
    END
  END vccd1.extra29
  PIN vccd1.extra30
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1624.020 -9.320 1627.020 430.000 ;
    END
  END vccd1.extra30
  PIN vccd1.extra31
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1444.020 -9.320 1447.020 430.000 ;
    END
  END vccd1.extra31
  PIN vccd1.extra32
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1264.020 -9.320 1267.020 430.000 ;
    END
  END vccd1.extra32
  PIN vccd1.extra33
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1084.020 -9.320 1087.020 430.000 ;
    END
  END vccd1.extra33
  PIN vccd1.extra34
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 904.020 -9.320 907.020 430.000 ;
    END
  END vccd1.extra34
  PIN vccd1.extra35
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 724.020 -9.320 727.020 430.000 ;
    END
  END vccd1.extra35
  PIN vccd1.extra36
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 544.020 -9.320 547.020 430.000 ;
    END
  END vccd1.extra36
  PIN vccd1.extra37
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 364.020 -9.320 367.020 430.000 ;
    END
  END vccd1.extra37
  PIN vccd1.extra38
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 3708.980 3529.900 3711.980 ;
    END
  END vccd1.extra38
  PIN vccd1.extra39
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3609.380 3534.600 3612.380 ;
    END
  END vccd1.extra39
  PIN vccd1.extra40
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3429.380 3534.600 3432.380 ;
    END
  END vccd1.extra40
  PIN vccd1.extra41
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3249.380 3534.600 3252.380 ;
    END
  END vccd1.extra41
  PIN vccd1.extra42
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3069.380 3534.600 3072.380 ;
    END
  END vccd1.extra42
  PIN vccd1.extra43
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2889.380 3534.600 2892.380 ;
    END
  END vccd1.extra43
  PIN vccd1.extra44
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2709.380 3534.600 2712.380 ;
    END
  END vccd1.extra44
  PIN vccd1.extra45
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2529.380 3534.600 2532.380 ;
    END
  END vccd1.extra45
  PIN vccd1.extra46
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2349.380 3534.600 2352.380 ;
    END
  END vccd1.extra46
  PIN vccd1.extra47
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2169.380 3534.600 2172.380 ;
    END
  END vccd1.extra47
  PIN vccd1.extra48
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1989.380 3534.600 1992.380 ;
    END
  END vccd1.extra48
  PIN vccd1.extra49
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1809.380 3534.600 1812.380 ;
    END
  END vccd1.extra49
  PIN vccd1.extra50
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1629.380 3534.600 1632.380 ;
    END
  END vccd1.extra50
  PIN vccd1.extra51
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1449.380 3534.600 1452.380 ;
    END
  END vccd1.extra51
  PIN vccd1.extra52
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1269.380 3534.600 1272.380 ;
    END
  END vccd1.extra52
  PIN vccd1.extra53
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1089.380 3534.600 1092.380 ;
    END
  END vccd1.extra53
  PIN vccd1.extra54
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 909.380 3534.600 912.380 ;
    END
  END vccd1.extra54
  PIN vccd1.extra55
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 729.380 3534.600 732.380 ;
    END
  END vccd1.extra55
  PIN vccd1.extra56
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 549.380 3534.600 552.380 ;
    END
  END vccd1.extra56
  PIN vccd1.extra57
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 369.380 3534.600 372.380 ;
    END
  END vccd1.extra57
  PIN vccd1.extra58
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 189.380 3534.600 192.380 ;
    END
  END vccd1.extra58
  PIN vccd1.extra59
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 9.380 3534.600 12.380 ;
    END
  END vccd1.extra59
  PIN vccd1.extra60
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 -4.620 3529.900 -1.620 ;
    END
  END vccd1.extra60
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3531.600 -9.320 3534.600 3716.680 ;
    END
  END vssd1
  PIN vssd1.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3334.020 -9.320 3337.020 3716.680 ;
    END
  END vssd1.extra1
  PIN vssd1.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3154.020 3669.800 3157.020 3716.680 ;
    END
  END vssd1.extra2
  PIN vssd1.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2974.020 3669.800 2977.020 3716.680 ;
    END
  END vssd1.extra3
  PIN vssd1.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2794.020 3669.800 2797.020 3716.680 ;
    END
  END vssd1.extra4
  PIN vssd1.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2614.020 3669.800 2617.020 3716.680 ;
    END
  END vssd1.extra5
  PIN vssd1.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2434.020 3669.800 2437.020 3716.680 ;
    END
  END vssd1.extra6
  PIN vssd1.extra7
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2254.020 3669.800 2257.020 3716.680 ;
    END
  END vssd1.extra7
  PIN vssd1.extra8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2074.020 3669.800 2077.020 3716.680 ;
    END
  END vssd1.extra8
  PIN vssd1.extra9
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1894.020 3669.800 1897.020 3716.680 ;
    END
  END vssd1.extra9
  PIN vssd1.extra10
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1714.020 3669.800 1717.020 3716.680 ;
    END
  END vssd1.extra10
  PIN vssd1.extra11
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1534.020 3669.800 1537.020 3716.680 ;
    END
  END vssd1.extra11
  PIN vssd1.extra12
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1354.020 3669.800 1357.020 3716.680 ;
    END
  END vssd1.extra12
  PIN vssd1.extra13
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1174.020 3669.800 1177.020 3716.680 ;
    END
  END vssd1.extra13
  PIN vssd1.extra14
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 994.020 3669.800 997.020 3716.680 ;
    END
  END vssd1.extra14
  PIN vssd1.extra15
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 814.020 3669.800 817.020 3716.680 ;
    END
  END vssd1.extra15
  PIN vssd1.extra16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 634.020 3669.800 637.020 3716.680 ;
    END
  END vssd1.extra16
  PIN vssd1.extra17
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 454.020 3669.800 457.020 3716.680 ;
    END
  END vssd1.extra17
  PIN vssd1.extra18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 274.020 -9.320 277.020 3716.680 ;
    END
  END vssd1.extra18
  PIN vssd1.extra19
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 94.020 -9.320 97.020 3716.680 ;
    END
  END vssd1.extra19
  PIN vssd1.extra20
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3716.680 ;
    END
  END vssd1.extra20
  PIN vssd1.extra21
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3154.020 -9.320 3157.020 430.000 ;
    END
  END vssd1.extra21
  PIN vssd1.extra22
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2974.020 -9.320 2977.020 430.000 ;
    END
  END vssd1.extra22
  PIN vssd1.extra23
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2794.020 -9.320 2797.020 430.000 ;
    END
  END vssd1.extra23
  PIN vssd1.extra24
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2614.020 -9.320 2617.020 430.000 ;
    END
  END vssd1.extra24
  PIN vssd1.extra25
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2434.020 -9.320 2437.020 430.000 ;
    END
  END vssd1.extra25
  PIN vssd1.extra26
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2254.020 -9.320 2257.020 430.000 ;
    END
  END vssd1.extra26
  PIN vssd1.extra27
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2074.020 -9.320 2077.020 430.000 ;
    END
  END vssd1.extra27
  PIN vssd1.extra28
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1894.020 -9.320 1897.020 430.000 ;
    END
  END vssd1.extra28
  PIN vssd1.extra29
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1714.020 -9.320 1717.020 430.000 ;
    END
  END vssd1.extra29
  PIN vssd1.extra30
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1534.020 -9.320 1537.020 430.000 ;
    END
  END vssd1.extra30
  PIN vssd1.extra31
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1354.020 -9.320 1357.020 430.000 ;
    END
  END vssd1.extra31
  PIN vssd1.extra32
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1174.020 -9.320 1177.020 430.000 ;
    END
  END vssd1.extra32
  PIN vssd1.extra33
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 994.020 -9.320 997.020 430.000 ;
    END
  END vssd1.extra33
  PIN vssd1.extra34
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 814.020 -9.320 817.020 430.000 ;
    END
  END vssd1.extra34
  PIN vssd1.extra35
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 634.020 -9.320 637.020 430.000 ;
    END
  END vssd1.extra35
  PIN vssd1.extra36
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 454.020 -9.320 457.020 430.000 ;
    END
  END vssd1.extra36
  PIN vssd1.extra37
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3713.680 3534.600 3716.680 ;
    END
  END vssd1.extra37
  PIN vssd1.extra38
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3519.380 3534.600 3522.380 ;
    END
  END vssd1.extra38
  PIN vssd1.extra39
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3339.380 3534.600 3342.380 ;
    END
  END vssd1.extra39
  PIN vssd1.extra40
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3159.380 3534.600 3162.380 ;
    END
  END vssd1.extra40
  PIN vssd1.extra41
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2979.380 3534.600 2982.380 ;
    END
  END vssd1.extra41
  PIN vssd1.extra42
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2799.380 3534.600 2802.380 ;
    END
  END vssd1.extra42
  PIN vssd1.extra43
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2619.380 3534.600 2622.380 ;
    END
  END vssd1.extra43
  PIN vssd1.extra44
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2439.380 3534.600 2442.380 ;
    END
  END vssd1.extra44
  PIN vssd1.extra45
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2259.380 3534.600 2262.380 ;
    END
  END vssd1.extra45
  PIN vssd1.extra46
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2079.380 3534.600 2082.380 ;
    END
  END vssd1.extra46
  PIN vssd1.extra47
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1899.380 3534.600 1902.380 ;
    END
  END vssd1.extra47
  PIN vssd1.extra48
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1719.380 3534.600 1722.380 ;
    END
  END vssd1.extra48
  PIN vssd1.extra49
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1539.380 3534.600 1542.380 ;
    END
  END vssd1.extra49
  PIN vssd1.extra50
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1359.380 3534.600 1362.380 ;
    END
  END vssd1.extra50
  PIN vssd1.extra51
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1179.380 3534.600 1182.380 ;
    END
  END vssd1.extra51
  PIN vssd1.extra52
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 999.380 3534.600 1002.380 ;
    END
  END vssd1.extra52
  PIN vssd1.extra53
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 819.380 3534.600 822.380 ;
    END
  END vssd1.extra53
  PIN vssd1.extra54
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 639.380 3534.600 642.380 ;
    END
  END vssd1.extra54
  PIN vssd1.extra55
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 459.380 3534.600 462.380 ;
    END
  END vssd1.extra55
  PIN vssd1.extra56
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 279.380 3534.600 282.380 ;
    END
  END vssd1.extra56
  PIN vssd1.extra57
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 99.380 3534.600 102.380 ;
    END
  END vssd1.extra57
  PIN vssd1.extra58
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 -9.320 3534.600 -6.320 ;
    END
  END vssd1.extra58
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3536.300 -14.020 3539.300 3721.380 ;
    END
  END vccd2
  PIN vccd2.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3721.380 ;
    END
  END vccd2.extra1
  PIN vccd2.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 3718.380 3539.300 3721.380 ;
    END
  END vccd2.extra2
  PIN vccd2.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 -14.020 3539.300 -11.020 ;
    END
  END vccd2.extra3
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3541.000 -18.720 3544.000 3726.080 ;
    END
  END vssd2
  PIN vssd2.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3726.080 ;
    END
  END vssd2.extra1
  PIN vssd2.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 3723.080 3544.000 3726.080 ;
    END
  END vssd2.extra2
  PIN vssd2.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 -18.720 3544.000 -15.720 ;
    END
  END vssd2.extra3
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3545.700 -23.420 3548.700 3730.780 ;
    END
  END vdda1
  PIN vdda1.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3730.780 ;
    END
  END vdda1.extra1
  PIN vdda1.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 3727.780 3548.700 3730.780 ;
    END
  END vdda1.extra2
  PIN vdda1.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 -23.420 3548.700 -20.420 ;
    END
  END vdda1.extra3
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3550.400 -28.120 3553.400 3735.480 ;
    END
  END vssa1
  PIN vssa1.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3735.480 ;
    END
  END vssa1.extra1
  PIN vssa1.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 3732.480 3553.400 3735.480 ;
    END
  END vssa1.extra2
  PIN vssa1.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 -28.120 3553.400 -25.120 ;
    END
  END vssa1.extra3
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3555.100 -32.820 3558.100 3740.180 ;
    END
  END vdda2
  PIN vdda2.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3740.180 ;
    END
  END vdda2.extra1
  PIN vdda2.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 3737.180 3558.100 3740.180 ;
    END
  END vdda2.extra2
  PIN vdda2.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 -32.820 3558.100 -29.820 ;
    END
  END vdda2.extra3
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3559.800 -37.520 3562.800 3744.880 ;
    END
  END vssa2
  PIN vssa2.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3744.880 ;
    END
  END vssa2.extra1
  PIN vssa2.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 3741.880 3562.800 3744.880 ;
    END
  END vssa2.extra2
  PIN vssa2.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 -37.520 3562.800 -34.520 ;
    END
  END vssa2.extra3
  OBS
      LAYER li1 ;
        RECT 337.785 14.025 3171.095 3661.375 ;
      LAYER met1 ;
        RECT 3.290 13.700 3516.170 3688.620 ;
      LAYER met2 ;
        RECT 3.320 3705.720 48.570 3706.000 ;
        RECT 49.410 3705.720 146.090 3706.000 ;
        RECT 146.930 3705.720 244.070 3706.000 ;
        RECT 244.910 3705.720 341.590 3706.000 ;
        RECT 342.430 3705.720 439.570 3706.000 ;
        RECT 440.410 3705.720 537.090 3706.000 ;
        RECT 537.930 3705.720 635.070 3706.000 ;
        RECT 635.910 3705.720 732.590 3706.000 ;
        RECT 733.430 3705.720 830.570 3706.000 ;
        RECT 831.410 3705.720 928.550 3706.000 ;
        RECT 929.390 3705.720 1026.070 3706.000 ;
        RECT 1026.910 3705.720 1124.050 3706.000 ;
        RECT 1124.890 3705.720 1221.570 3706.000 ;
        RECT 1222.410 3705.720 1319.550 3706.000 ;
        RECT 1320.390 3705.720 1417.070 3706.000 ;
        RECT 1417.910 3705.720 1515.050 3706.000 ;
        RECT 1515.890 3705.720 1612.570 3706.000 ;
        RECT 1613.410 3705.720 1710.550 3706.000 ;
        RECT 1711.390 3705.720 1808.530 3706.000 ;
        RECT 1809.370 3705.720 1906.050 3706.000 ;
        RECT 1906.890 3705.720 2004.030 3706.000 ;
        RECT 2004.870 3705.720 2101.550 3706.000 ;
        RECT 2102.390 3705.720 2199.530 3706.000 ;
        RECT 2200.370 3705.720 2297.050 3706.000 ;
        RECT 2297.890 3705.720 2395.030 3706.000 ;
        RECT 2395.870 3705.720 2492.550 3706.000 ;
        RECT 2493.390 3705.720 2590.530 3706.000 ;
        RECT 2591.370 3705.720 2688.510 3706.000 ;
        RECT 2689.350 3705.720 2786.030 3706.000 ;
        RECT 2786.870 3705.720 2884.010 3706.000 ;
        RECT 2884.850 3705.720 2981.530 3706.000 ;
        RECT 2982.370 3705.720 3079.510 3706.000 ;
        RECT 3080.350 3705.720 3177.030 3706.000 ;
        RECT 3177.870 3705.720 3275.010 3706.000 ;
        RECT 3275.850 3705.720 3372.530 3706.000 ;
        RECT 3373.370 3705.720 3470.510 3706.000 ;
        RECT 3471.350 3705.720 3516.140 3706.000 ;
        RECT 3.320 4.280 3516.140 3705.720 ;
        RECT 3.870 4.000 9.930 4.280 ;
        RECT 10.770 4.000 16.830 4.280 ;
        RECT 17.670 4.000 24.190 4.280 ;
        RECT 25.030 4.000 31.090 4.280 ;
        RECT 31.930 4.000 38.450 4.280 ;
        RECT 39.290 4.000 45.350 4.280 ;
        RECT 46.190 4.000 52.710 4.280 ;
        RECT 53.550 4.000 59.610 4.280 ;
        RECT 60.450 4.000 66.970 4.280 ;
        RECT 67.810 4.000 73.870 4.280 ;
        RECT 74.710 4.000 81.230 4.280 ;
        RECT 82.070 4.000 88.130 4.280 ;
        RECT 88.970 4.000 95.490 4.280 ;
        RECT 96.330 4.000 102.390 4.280 ;
        RECT 103.230 4.000 109.750 4.280 ;
        RECT 110.590 4.000 116.650 4.280 ;
        RECT 117.490 4.000 124.010 4.280 ;
        RECT 124.850 4.000 130.910 4.280 ;
        RECT 131.750 4.000 138.270 4.280 ;
        RECT 139.110 4.000 145.170 4.280 ;
        RECT 146.010 4.000 152.530 4.280 ;
        RECT 153.370 4.000 159.430 4.280 ;
        RECT 160.270 4.000 166.790 4.280 ;
        RECT 167.630 4.000 173.690 4.280 ;
        RECT 174.530 4.000 181.050 4.280 ;
        RECT 181.890 4.000 187.950 4.280 ;
        RECT 188.790 4.000 195.310 4.280 ;
        RECT 196.150 4.000 202.210 4.280 ;
        RECT 203.050 4.000 209.570 4.280 ;
        RECT 210.410 4.000 216.470 4.280 ;
        RECT 217.310 4.000 223.830 4.280 ;
        RECT 224.670 4.000 230.730 4.280 ;
        RECT 231.570 4.000 238.090 4.280 ;
        RECT 238.930 4.000 244.990 4.280 ;
        RECT 245.830 4.000 252.350 4.280 ;
        RECT 253.190 4.000 259.250 4.280 ;
        RECT 260.090 4.000 266.610 4.280 ;
        RECT 267.450 4.000 273.510 4.280 ;
        RECT 274.350 4.000 280.870 4.280 ;
        RECT 281.710 4.000 287.770 4.280 ;
        RECT 288.610 4.000 295.130 4.280 ;
        RECT 295.970 4.000 302.030 4.280 ;
        RECT 302.870 4.000 309.390 4.280 ;
        RECT 310.230 4.000 316.290 4.280 ;
        RECT 317.130 4.000 323.650 4.280 ;
        RECT 324.490 4.000 330.550 4.280 ;
        RECT 331.390 4.000 337.910 4.280 ;
        RECT 338.750 4.000 344.810 4.280 ;
        RECT 345.650 4.000 352.170 4.280 ;
        RECT 353.010 4.000 359.070 4.280 ;
        RECT 359.910 4.000 365.970 4.280 ;
        RECT 366.810 4.000 373.330 4.280 ;
        RECT 374.170 4.000 380.230 4.280 ;
        RECT 381.070 4.000 387.590 4.280 ;
        RECT 388.430 4.000 394.490 4.280 ;
        RECT 395.330 4.000 401.850 4.280 ;
        RECT 402.690 4.000 408.750 4.280 ;
        RECT 409.590 4.000 416.110 4.280 ;
        RECT 416.950 4.000 423.010 4.280 ;
        RECT 423.850 4.000 430.370 4.280 ;
        RECT 431.210 4.000 437.270 4.280 ;
        RECT 438.110 4.000 444.630 4.280 ;
        RECT 445.470 4.000 451.530 4.280 ;
        RECT 452.370 4.000 458.890 4.280 ;
        RECT 459.730 4.000 465.790 4.280 ;
        RECT 466.630 4.000 473.150 4.280 ;
        RECT 473.990 4.000 480.050 4.280 ;
        RECT 480.890 4.000 487.410 4.280 ;
        RECT 488.250 4.000 494.310 4.280 ;
        RECT 495.150 4.000 501.670 4.280 ;
        RECT 502.510 4.000 508.570 4.280 ;
        RECT 509.410 4.000 515.930 4.280 ;
        RECT 516.770 4.000 522.830 4.280 ;
        RECT 523.670 4.000 530.190 4.280 ;
        RECT 531.030 4.000 537.090 4.280 ;
        RECT 537.930 4.000 544.450 4.280 ;
        RECT 545.290 4.000 551.350 4.280 ;
        RECT 552.190 4.000 558.710 4.280 ;
        RECT 559.550 4.000 565.610 4.280 ;
        RECT 566.450 4.000 572.970 4.280 ;
        RECT 573.810 4.000 579.870 4.280 ;
        RECT 580.710 4.000 587.230 4.280 ;
        RECT 588.070 4.000 594.130 4.280 ;
        RECT 594.970 4.000 601.490 4.280 ;
        RECT 602.330 4.000 608.390 4.280 ;
        RECT 609.230 4.000 615.750 4.280 ;
        RECT 616.590 4.000 622.650 4.280 ;
        RECT 623.490 4.000 630.010 4.280 ;
        RECT 630.850 4.000 636.910 4.280 ;
        RECT 637.750 4.000 644.270 4.280 ;
        RECT 645.110 4.000 651.170 4.280 ;
        RECT 652.010 4.000 658.530 4.280 ;
        RECT 659.370 4.000 665.430 4.280 ;
        RECT 666.270 4.000 672.790 4.280 ;
        RECT 673.630 4.000 679.690 4.280 ;
        RECT 680.530 4.000 687.050 4.280 ;
        RECT 687.890 4.000 693.950 4.280 ;
        RECT 694.790 4.000 701.310 4.280 ;
        RECT 702.150 4.000 708.210 4.280 ;
        RECT 709.050 4.000 715.110 4.280 ;
        RECT 715.950 4.000 722.470 4.280 ;
        RECT 723.310 4.000 729.370 4.280 ;
        RECT 730.210 4.000 736.730 4.280 ;
        RECT 737.570 4.000 743.630 4.280 ;
        RECT 744.470 4.000 750.990 4.280 ;
        RECT 751.830 4.000 757.890 4.280 ;
        RECT 758.730 4.000 765.250 4.280 ;
        RECT 766.090 4.000 772.150 4.280 ;
        RECT 772.990 4.000 779.510 4.280 ;
        RECT 780.350 4.000 786.410 4.280 ;
        RECT 787.250 4.000 793.770 4.280 ;
        RECT 794.610 4.000 800.670 4.280 ;
        RECT 801.510 4.000 808.030 4.280 ;
        RECT 808.870 4.000 814.930 4.280 ;
        RECT 815.770 4.000 822.290 4.280 ;
        RECT 823.130 4.000 829.190 4.280 ;
        RECT 830.030 4.000 836.550 4.280 ;
        RECT 837.390 4.000 843.450 4.280 ;
        RECT 844.290 4.000 850.810 4.280 ;
        RECT 851.650 4.000 857.710 4.280 ;
        RECT 858.550 4.000 865.070 4.280 ;
        RECT 865.910 4.000 871.970 4.280 ;
        RECT 872.810 4.000 879.330 4.280 ;
        RECT 880.170 4.000 886.230 4.280 ;
        RECT 887.070 4.000 893.590 4.280 ;
        RECT 894.430 4.000 900.490 4.280 ;
        RECT 901.330 4.000 907.850 4.280 ;
        RECT 908.690 4.000 914.750 4.280 ;
        RECT 915.590 4.000 922.110 4.280 ;
        RECT 922.950 4.000 929.010 4.280 ;
        RECT 929.850 4.000 936.370 4.280 ;
        RECT 937.210 4.000 943.270 4.280 ;
        RECT 944.110 4.000 950.630 4.280 ;
        RECT 951.470 4.000 957.530 4.280 ;
        RECT 958.370 4.000 964.890 4.280 ;
        RECT 965.730 4.000 971.790 4.280 ;
        RECT 972.630 4.000 979.150 4.280 ;
        RECT 979.990 4.000 986.050 4.280 ;
        RECT 986.890 4.000 993.410 4.280 ;
        RECT 994.250 4.000 1000.310 4.280 ;
        RECT 1001.150 4.000 1007.670 4.280 ;
        RECT 1008.510 4.000 1014.570 4.280 ;
        RECT 1015.410 4.000 1021.930 4.280 ;
        RECT 1022.770 4.000 1028.830 4.280 ;
        RECT 1029.670 4.000 1036.190 4.280 ;
        RECT 1037.030 4.000 1043.090 4.280 ;
        RECT 1043.930 4.000 1050.450 4.280 ;
        RECT 1051.290 4.000 1057.350 4.280 ;
        RECT 1058.190 4.000 1064.250 4.280 ;
        RECT 1065.090 4.000 1071.610 4.280 ;
        RECT 1072.450 4.000 1078.510 4.280 ;
        RECT 1079.350 4.000 1085.870 4.280 ;
        RECT 1086.710 4.000 1092.770 4.280 ;
        RECT 1093.610 4.000 1100.130 4.280 ;
        RECT 1100.970 4.000 1107.030 4.280 ;
        RECT 1107.870 4.000 1114.390 4.280 ;
        RECT 1115.230 4.000 1121.290 4.280 ;
        RECT 1122.130 4.000 1128.650 4.280 ;
        RECT 1129.490 4.000 1135.550 4.280 ;
        RECT 1136.390 4.000 1142.910 4.280 ;
        RECT 1143.750 4.000 1149.810 4.280 ;
        RECT 1150.650 4.000 1157.170 4.280 ;
        RECT 1158.010 4.000 1164.070 4.280 ;
        RECT 1164.910 4.000 1171.430 4.280 ;
        RECT 1172.270 4.000 1178.330 4.280 ;
        RECT 1179.170 4.000 1185.690 4.280 ;
        RECT 1186.530 4.000 1192.590 4.280 ;
        RECT 1193.430 4.000 1199.950 4.280 ;
        RECT 1200.790 4.000 1206.850 4.280 ;
        RECT 1207.690 4.000 1214.210 4.280 ;
        RECT 1215.050 4.000 1221.110 4.280 ;
        RECT 1221.950 4.000 1228.470 4.280 ;
        RECT 1229.310 4.000 1235.370 4.280 ;
        RECT 1236.210 4.000 1242.730 4.280 ;
        RECT 1243.570 4.000 1249.630 4.280 ;
        RECT 1250.470 4.000 1256.990 4.280 ;
        RECT 1257.830 4.000 1263.890 4.280 ;
        RECT 1264.730 4.000 1271.250 4.280 ;
        RECT 1272.090 4.000 1278.150 4.280 ;
        RECT 1278.990 4.000 1285.510 4.280 ;
        RECT 1286.350 4.000 1292.410 4.280 ;
        RECT 1293.250 4.000 1299.770 4.280 ;
        RECT 1300.610 4.000 1306.670 4.280 ;
        RECT 1307.510 4.000 1314.030 4.280 ;
        RECT 1314.870 4.000 1320.930 4.280 ;
        RECT 1321.770 4.000 1328.290 4.280 ;
        RECT 1329.130 4.000 1335.190 4.280 ;
        RECT 1336.030 4.000 1342.550 4.280 ;
        RECT 1343.390 4.000 1349.450 4.280 ;
        RECT 1350.290 4.000 1356.810 4.280 ;
        RECT 1357.650 4.000 1363.710 4.280 ;
        RECT 1364.550 4.000 1371.070 4.280 ;
        RECT 1371.910 4.000 1377.970 4.280 ;
        RECT 1378.810 4.000 1385.330 4.280 ;
        RECT 1386.170 4.000 1392.230 4.280 ;
        RECT 1393.070 4.000 1399.590 4.280 ;
        RECT 1400.430 4.000 1406.490 4.280 ;
        RECT 1407.330 4.000 1413.390 4.280 ;
        RECT 1414.230 4.000 1420.750 4.280 ;
        RECT 1421.590 4.000 1427.650 4.280 ;
        RECT 1428.490 4.000 1435.010 4.280 ;
        RECT 1435.850 4.000 1441.910 4.280 ;
        RECT 1442.750 4.000 1449.270 4.280 ;
        RECT 1450.110 4.000 1456.170 4.280 ;
        RECT 1457.010 4.000 1463.530 4.280 ;
        RECT 1464.370 4.000 1470.430 4.280 ;
        RECT 1471.270 4.000 1477.790 4.280 ;
        RECT 1478.630 4.000 1484.690 4.280 ;
        RECT 1485.530 4.000 1492.050 4.280 ;
        RECT 1492.890 4.000 1498.950 4.280 ;
        RECT 1499.790 4.000 1506.310 4.280 ;
        RECT 1507.150 4.000 1513.210 4.280 ;
        RECT 1514.050 4.000 1520.570 4.280 ;
        RECT 1521.410 4.000 1527.470 4.280 ;
        RECT 1528.310 4.000 1534.830 4.280 ;
        RECT 1535.670 4.000 1541.730 4.280 ;
        RECT 1542.570 4.000 1549.090 4.280 ;
        RECT 1549.930 4.000 1555.990 4.280 ;
        RECT 1556.830 4.000 1563.350 4.280 ;
        RECT 1564.190 4.000 1570.250 4.280 ;
        RECT 1571.090 4.000 1577.610 4.280 ;
        RECT 1578.450 4.000 1584.510 4.280 ;
        RECT 1585.350 4.000 1591.870 4.280 ;
        RECT 1592.710 4.000 1598.770 4.280 ;
        RECT 1599.610 4.000 1606.130 4.280 ;
        RECT 1606.970 4.000 1613.030 4.280 ;
        RECT 1613.870 4.000 1620.390 4.280 ;
        RECT 1621.230 4.000 1627.290 4.280 ;
        RECT 1628.130 4.000 1634.650 4.280 ;
        RECT 1635.490 4.000 1641.550 4.280 ;
        RECT 1642.390 4.000 1648.910 4.280 ;
        RECT 1649.750 4.000 1655.810 4.280 ;
        RECT 1656.650 4.000 1663.170 4.280 ;
        RECT 1664.010 4.000 1670.070 4.280 ;
        RECT 1670.910 4.000 1677.430 4.280 ;
        RECT 1678.270 4.000 1684.330 4.280 ;
        RECT 1685.170 4.000 1691.690 4.280 ;
        RECT 1692.530 4.000 1698.590 4.280 ;
        RECT 1699.430 4.000 1705.950 4.280 ;
        RECT 1706.790 4.000 1712.850 4.280 ;
        RECT 1713.690 4.000 1720.210 4.280 ;
        RECT 1721.050 4.000 1727.110 4.280 ;
        RECT 1727.950 4.000 1734.470 4.280 ;
        RECT 1735.310 4.000 1741.370 4.280 ;
        RECT 1742.210 4.000 1748.730 4.280 ;
        RECT 1749.570 4.000 1755.630 4.280 ;
        RECT 1756.470 4.000 1762.990 4.280 ;
        RECT 1763.830 4.000 1769.890 4.280 ;
        RECT 1770.730 4.000 1776.790 4.280 ;
        RECT 1777.630 4.000 1784.150 4.280 ;
        RECT 1784.990 4.000 1791.050 4.280 ;
        RECT 1791.890 4.000 1798.410 4.280 ;
        RECT 1799.250 4.000 1805.310 4.280 ;
        RECT 1806.150 4.000 1812.670 4.280 ;
        RECT 1813.510 4.000 1819.570 4.280 ;
        RECT 1820.410 4.000 1826.930 4.280 ;
        RECT 1827.770 4.000 1833.830 4.280 ;
        RECT 1834.670 4.000 1841.190 4.280 ;
        RECT 1842.030 4.000 1848.090 4.280 ;
        RECT 1848.930 4.000 1855.450 4.280 ;
        RECT 1856.290 4.000 1862.350 4.280 ;
        RECT 1863.190 4.000 1869.710 4.280 ;
        RECT 1870.550 4.000 1876.610 4.280 ;
        RECT 1877.450 4.000 1883.970 4.280 ;
        RECT 1884.810 4.000 1890.870 4.280 ;
        RECT 1891.710 4.000 1898.230 4.280 ;
        RECT 1899.070 4.000 1905.130 4.280 ;
        RECT 1905.970 4.000 1912.490 4.280 ;
        RECT 1913.330 4.000 1919.390 4.280 ;
        RECT 1920.230 4.000 1926.750 4.280 ;
        RECT 1927.590 4.000 1933.650 4.280 ;
        RECT 1934.490 4.000 1941.010 4.280 ;
        RECT 1941.850 4.000 1947.910 4.280 ;
        RECT 1948.750 4.000 1955.270 4.280 ;
        RECT 1956.110 4.000 1962.170 4.280 ;
        RECT 1963.010 4.000 1969.530 4.280 ;
        RECT 1970.370 4.000 1976.430 4.280 ;
        RECT 1977.270 4.000 1983.790 4.280 ;
        RECT 1984.630 4.000 1990.690 4.280 ;
        RECT 1991.530 4.000 1998.050 4.280 ;
        RECT 1998.890 4.000 2004.950 4.280 ;
        RECT 2005.790 4.000 2012.310 4.280 ;
        RECT 2013.150 4.000 2019.210 4.280 ;
        RECT 2020.050 4.000 2026.570 4.280 ;
        RECT 2027.410 4.000 2033.470 4.280 ;
        RECT 2034.310 4.000 2040.830 4.280 ;
        RECT 2041.670 4.000 2047.730 4.280 ;
        RECT 2048.570 4.000 2055.090 4.280 ;
        RECT 2055.930 4.000 2061.990 4.280 ;
        RECT 2062.830 4.000 2069.350 4.280 ;
        RECT 2070.190 4.000 2076.250 4.280 ;
        RECT 2077.090 4.000 2083.610 4.280 ;
        RECT 2084.450 4.000 2090.510 4.280 ;
        RECT 2091.350 4.000 2097.870 4.280 ;
        RECT 2098.710 4.000 2104.770 4.280 ;
        RECT 2105.610 4.000 2112.130 4.280 ;
        RECT 2112.970 4.000 2119.030 4.280 ;
        RECT 2119.870 4.000 2125.930 4.280 ;
        RECT 2126.770 4.000 2133.290 4.280 ;
        RECT 2134.130 4.000 2140.190 4.280 ;
        RECT 2141.030 4.000 2147.550 4.280 ;
        RECT 2148.390 4.000 2154.450 4.280 ;
        RECT 2155.290 4.000 2161.810 4.280 ;
        RECT 2162.650 4.000 2168.710 4.280 ;
        RECT 2169.550 4.000 2176.070 4.280 ;
        RECT 2176.910 4.000 2182.970 4.280 ;
        RECT 2183.810 4.000 2190.330 4.280 ;
        RECT 2191.170 4.000 2197.230 4.280 ;
        RECT 2198.070 4.000 2204.590 4.280 ;
        RECT 2205.430 4.000 2211.490 4.280 ;
        RECT 2212.330 4.000 2218.850 4.280 ;
        RECT 2219.690 4.000 2225.750 4.280 ;
        RECT 2226.590 4.000 2233.110 4.280 ;
        RECT 2233.950 4.000 2240.010 4.280 ;
        RECT 2240.850 4.000 2247.370 4.280 ;
        RECT 2248.210 4.000 2254.270 4.280 ;
        RECT 2255.110 4.000 2261.630 4.280 ;
        RECT 2262.470 4.000 2268.530 4.280 ;
        RECT 2269.370 4.000 2275.890 4.280 ;
        RECT 2276.730 4.000 2282.790 4.280 ;
        RECT 2283.630 4.000 2290.150 4.280 ;
        RECT 2290.990 4.000 2297.050 4.280 ;
        RECT 2297.890 4.000 2304.410 4.280 ;
        RECT 2305.250 4.000 2311.310 4.280 ;
        RECT 2312.150 4.000 2318.670 4.280 ;
        RECT 2319.510 4.000 2325.570 4.280 ;
        RECT 2326.410 4.000 2332.930 4.280 ;
        RECT 2333.770 4.000 2339.830 4.280 ;
        RECT 2340.670 4.000 2347.190 4.280 ;
        RECT 2348.030 4.000 2354.090 4.280 ;
        RECT 2354.930 4.000 2361.450 4.280 ;
        RECT 2362.290 4.000 2368.350 4.280 ;
        RECT 2369.190 4.000 2375.710 4.280 ;
        RECT 2376.550 4.000 2382.610 4.280 ;
        RECT 2383.450 4.000 2389.970 4.280 ;
        RECT 2390.810 4.000 2396.870 4.280 ;
        RECT 2397.710 4.000 2404.230 4.280 ;
        RECT 2405.070 4.000 2411.130 4.280 ;
        RECT 2411.970 4.000 2418.490 4.280 ;
        RECT 2419.330 4.000 2425.390 4.280 ;
        RECT 2426.230 4.000 2432.750 4.280 ;
        RECT 2433.590 4.000 2439.650 4.280 ;
        RECT 2440.490 4.000 2447.010 4.280 ;
        RECT 2447.850 4.000 2453.910 4.280 ;
        RECT 2454.750 4.000 2461.270 4.280 ;
        RECT 2462.110 4.000 2468.170 4.280 ;
        RECT 2469.010 4.000 2475.070 4.280 ;
        RECT 2475.910 4.000 2482.430 4.280 ;
        RECT 2483.270 4.000 2489.330 4.280 ;
        RECT 2490.170 4.000 2496.690 4.280 ;
        RECT 2497.530 4.000 2503.590 4.280 ;
        RECT 2504.430 4.000 2510.950 4.280 ;
        RECT 2511.790 4.000 2517.850 4.280 ;
        RECT 2518.690 4.000 2525.210 4.280 ;
        RECT 2526.050 4.000 2532.110 4.280 ;
        RECT 2532.950 4.000 2539.470 4.280 ;
        RECT 2540.310 4.000 2546.370 4.280 ;
        RECT 2547.210 4.000 2553.730 4.280 ;
        RECT 2554.570 4.000 2560.630 4.280 ;
        RECT 2561.470 4.000 2567.990 4.280 ;
        RECT 2568.830 4.000 2574.890 4.280 ;
        RECT 2575.730 4.000 2582.250 4.280 ;
        RECT 2583.090 4.000 2589.150 4.280 ;
        RECT 2589.990 4.000 2596.510 4.280 ;
        RECT 2597.350 4.000 2603.410 4.280 ;
        RECT 2604.250 4.000 2610.770 4.280 ;
        RECT 2611.610 4.000 2617.670 4.280 ;
        RECT 2618.510 4.000 2625.030 4.280 ;
        RECT 2625.870 4.000 2631.930 4.280 ;
        RECT 2632.770 4.000 2639.290 4.280 ;
        RECT 2640.130 4.000 2646.190 4.280 ;
        RECT 2647.030 4.000 2653.550 4.280 ;
        RECT 2654.390 4.000 2660.450 4.280 ;
        RECT 2661.290 4.000 2667.810 4.280 ;
        RECT 2668.650 4.000 2674.710 4.280 ;
        RECT 2675.550 4.000 2682.070 4.280 ;
        RECT 2682.910 4.000 2688.970 4.280 ;
        RECT 2689.810 4.000 2696.330 4.280 ;
        RECT 2697.170 4.000 2703.230 4.280 ;
        RECT 2704.070 4.000 2710.590 4.280 ;
        RECT 2711.430 4.000 2717.490 4.280 ;
        RECT 2718.330 4.000 2724.850 4.280 ;
        RECT 2725.690 4.000 2731.750 4.280 ;
        RECT 2732.590 4.000 2739.110 4.280 ;
        RECT 2739.950 4.000 2746.010 4.280 ;
        RECT 2746.850 4.000 2753.370 4.280 ;
        RECT 2754.210 4.000 2760.270 4.280 ;
        RECT 2761.110 4.000 2767.630 4.280 ;
        RECT 2768.470 4.000 2774.530 4.280 ;
        RECT 2775.370 4.000 2781.890 4.280 ;
        RECT 2782.730 4.000 2788.790 4.280 ;
        RECT 2789.630 4.000 2796.150 4.280 ;
        RECT 2796.990 4.000 2803.050 4.280 ;
        RECT 2803.890 4.000 2810.410 4.280 ;
        RECT 2811.250 4.000 2817.310 4.280 ;
        RECT 2818.150 4.000 2824.210 4.280 ;
        RECT 2825.050 4.000 2831.570 4.280 ;
        RECT 2832.410 4.000 2838.470 4.280 ;
        RECT 2839.310 4.000 2845.830 4.280 ;
        RECT 2846.670 4.000 2852.730 4.280 ;
        RECT 2853.570 4.000 2860.090 4.280 ;
        RECT 2860.930 4.000 2866.990 4.280 ;
        RECT 2867.830 4.000 2874.350 4.280 ;
        RECT 2875.190 4.000 2881.250 4.280 ;
        RECT 2882.090 4.000 2888.610 4.280 ;
        RECT 2889.450 4.000 2895.510 4.280 ;
        RECT 2896.350 4.000 2902.870 4.280 ;
        RECT 2903.710 4.000 2909.770 4.280 ;
        RECT 2910.610 4.000 2917.130 4.280 ;
        RECT 2917.970 4.000 2924.030 4.280 ;
        RECT 2924.870 4.000 2931.390 4.280 ;
        RECT 2932.230 4.000 2938.290 4.280 ;
        RECT 2939.130 4.000 2945.650 4.280 ;
        RECT 2946.490 4.000 2952.550 4.280 ;
        RECT 2953.390 4.000 2959.910 4.280 ;
        RECT 2960.750 4.000 2966.810 4.280 ;
        RECT 2967.650 4.000 2974.170 4.280 ;
        RECT 2975.010 4.000 2981.070 4.280 ;
        RECT 2981.910 4.000 2988.430 4.280 ;
        RECT 2989.270 4.000 2995.330 4.280 ;
        RECT 2996.170 4.000 3002.690 4.280 ;
        RECT 3003.530 4.000 3009.590 4.280 ;
        RECT 3010.430 4.000 3016.950 4.280 ;
        RECT 3017.790 4.000 3023.850 4.280 ;
        RECT 3024.690 4.000 3031.210 4.280 ;
        RECT 3032.050 4.000 3038.110 4.280 ;
        RECT 3038.950 4.000 3045.470 4.280 ;
        RECT 3046.310 4.000 3052.370 4.280 ;
        RECT 3053.210 4.000 3059.730 4.280 ;
        RECT 3060.570 4.000 3066.630 4.280 ;
        RECT 3067.470 4.000 3073.990 4.280 ;
        RECT 3074.830 4.000 3080.890 4.280 ;
        RECT 3081.730 4.000 3088.250 4.280 ;
        RECT 3089.090 4.000 3095.150 4.280 ;
        RECT 3095.990 4.000 3102.510 4.280 ;
        RECT 3103.350 4.000 3109.410 4.280 ;
        RECT 3110.250 4.000 3116.770 4.280 ;
        RECT 3117.610 4.000 3123.670 4.280 ;
        RECT 3124.510 4.000 3131.030 4.280 ;
        RECT 3131.870 4.000 3137.930 4.280 ;
        RECT 3138.770 4.000 3145.290 4.280 ;
        RECT 3146.130 4.000 3152.190 4.280 ;
        RECT 3153.030 4.000 3159.550 4.280 ;
        RECT 3160.390 4.000 3166.450 4.280 ;
        RECT 3167.290 4.000 3173.350 4.280 ;
        RECT 3174.190 4.000 3180.710 4.280 ;
        RECT 3181.550 4.000 3187.610 4.280 ;
        RECT 3188.450 4.000 3194.970 4.280 ;
        RECT 3195.810 4.000 3201.870 4.280 ;
        RECT 3202.710 4.000 3209.230 4.280 ;
        RECT 3210.070 4.000 3216.130 4.280 ;
        RECT 3216.970 4.000 3223.490 4.280 ;
        RECT 3224.330 4.000 3230.390 4.280 ;
        RECT 3231.230 4.000 3237.750 4.280 ;
        RECT 3238.590 4.000 3244.650 4.280 ;
        RECT 3245.490 4.000 3252.010 4.280 ;
        RECT 3252.850 4.000 3258.910 4.280 ;
        RECT 3259.750 4.000 3266.270 4.280 ;
        RECT 3267.110 4.000 3273.170 4.280 ;
        RECT 3274.010 4.000 3280.530 4.280 ;
        RECT 3281.370 4.000 3287.430 4.280 ;
        RECT 3288.270 4.000 3294.790 4.280 ;
        RECT 3295.630 4.000 3301.690 4.280 ;
        RECT 3302.530 4.000 3309.050 4.280 ;
        RECT 3309.890 4.000 3315.950 4.280 ;
        RECT 3316.790 4.000 3323.310 4.280 ;
        RECT 3324.150 4.000 3330.210 4.280 ;
        RECT 3331.050 4.000 3337.570 4.280 ;
        RECT 3338.410 4.000 3344.470 4.280 ;
        RECT 3345.310 4.000 3351.830 4.280 ;
        RECT 3352.670 4.000 3358.730 4.280 ;
        RECT 3359.570 4.000 3366.090 4.280 ;
        RECT 3366.930 4.000 3372.990 4.280 ;
        RECT 3373.830 4.000 3380.350 4.280 ;
        RECT 3381.190 4.000 3387.250 4.280 ;
        RECT 3388.090 4.000 3394.610 4.280 ;
        RECT 3395.450 4.000 3401.510 4.280 ;
        RECT 3402.350 4.000 3408.870 4.280 ;
        RECT 3409.710 4.000 3415.770 4.280 ;
        RECT 3416.610 4.000 3423.130 4.280 ;
        RECT 3423.970 4.000 3430.030 4.280 ;
        RECT 3430.870 4.000 3437.390 4.280 ;
        RECT 3438.230 4.000 3444.290 4.280 ;
        RECT 3445.130 4.000 3451.650 4.280 ;
        RECT 3452.490 4.000 3458.550 4.280 ;
        RECT 3459.390 4.000 3465.910 4.280 ;
        RECT 3466.750 4.000 3472.810 4.280 ;
        RECT 3473.650 4.000 3480.170 4.280 ;
        RECT 3481.010 4.000 3487.070 4.280 ;
        RECT 3487.910 4.000 3494.430 4.280 ;
        RECT 3495.270 4.000 3501.330 4.280 ;
        RECT 3502.170 4.000 3508.690 4.280 ;
        RECT 3509.530 4.000 3515.590 4.280 ;
      LAYER met3 ;
        RECT 4.400 3674.360 3515.600 3675.225 ;
        RECT 4.000 3607.080 3516.000 3674.360 ;
        RECT 4.400 3605.720 3516.000 3607.080 ;
        RECT 4.400 3605.680 3515.600 3605.720 ;
        RECT 4.000 3604.320 3515.600 3605.680 ;
        RECT 4.000 3538.400 3516.000 3604.320 ;
        RECT 4.400 3537.000 3516.000 3538.400 ;
        RECT 4.000 3535.680 3516.000 3537.000 ;
        RECT 4.000 3534.280 3515.600 3535.680 ;
        RECT 4.000 3469.720 3516.000 3534.280 ;
        RECT 4.400 3468.320 3516.000 3469.720 ;
        RECT 4.000 3465.640 3516.000 3468.320 ;
        RECT 4.000 3464.240 3515.600 3465.640 ;
        RECT 4.000 3401.040 3516.000 3464.240 ;
        RECT 4.400 3399.640 3516.000 3401.040 ;
        RECT 4.000 3395.600 3516.000 3399.640 ;
        RECT 4.000 3394.200 3515.600 3395.600 ;
        RECT 4.000 3332.360 3516.000 3394.200 ;
        RECT 4.400 3330.960 3516.000 3332.360 ;
        RECT 4.000 3325.560 3516.000 3330.960 ;
        RECT 4.000 3324.160 3515.600 3325.560 ;
        RECT 4.000 3263.680 3516.000 3324.160 ;
        RECT 4.400 3262.280 3516.000 3263.680 ;
        RECT 4.000 3255.520 3516.000 3262.280 ;
        RECT 4.000 3254.120 3515.600 3255.520 ;
        RECT 4.000 3195.000 3516.000 3254.120 ;
        RECT 4.400 3193.600 3516.000 3195.000 ;
        RECT 4.000 3185.480 3516.000 3193.600 ;
        RECT 4.000 3184.080 3515.600 3185.480 ;
        RECT 4.000 3126.320 3516.000 3184.080 ;
        RECT 4.400 3124.920 3516.000 3126.320 ;
        RECT 4.000 3115.440 3516.000 3124.920 ;
        RECT 4.000 3114.040 3515.600 3115.440 ;
        RECT 4.000 3057.640 3516.000 3114.040 ;
        RECT 4.400 3056.240 3516.000 3057.640 ;
        RECT 4.000 3045.400 3516.000 3056.240 ;
        RECT 4.000 3044.000 3515.600 3045.400 ;
        RECT 4.000 2988.960 3516.000 3044.000 ;
        RECT 4.400 2987.560 3516.000 2988.960 ;
        RECT 4.000 2975.360 3516.000 2987.560 ;
        RECT 4.000 2973.960 3515.600 2975.360 ;
        RECT 4.000 2920.280 3516.000 2973.960 ;
        RECT 4.400 2918.880 3516.000 2920.280 ;
        RECT 4.000 2905.320 3516.000 2918.880 ;
        RECT 4.000 2903.920 3515.600 2905.320 ;
        RECT 4.000 2851.600 3516.000 2903.920 ;
        RECT 4.400 2850.200 3516.000 2851.600 ;
        RECT 4.000 2835.280 3516.000 2850.200 ;
        RECT 4.000 2833.880 3515.600 2835.280 ;
        RECT 4.000 2782.920 3516.000 2833.880 ;
        RECT 4.400 2781.520 3516.000 2782.920 ;
        RECT 4.000 2765.240 3516.000 2781.520 ;
        RECT 4.000 2763.840 3515.600 2765.240 ;
        RECT 4.000 2714.240 3516.000 2763.840 ;
        RECT 4.400 2712.840 3516.000 2714.240 ;
        RECT 4.000 2695.200 3516.000 2712.840 ;
        RECT 4.000 2693.800 3515.600 2695.200 ;
        RECT 4.000 2645.560 3516.000 2693.800 ;
        RECT 4.400 2644.160 3516.000 2645.560 ;
        RECT 4.000 2625.160 3516.000 2644.160 ;
        RECT 4.000 2623.760 3515.600 2625.160 ;
        RECT 4.000 2576.880 3516.000 2623.760 ;
        RECT 4.400 2575.480 3516.000 2576.880 ;
        RECT 4.000 2555.120 3516.000 2575.480 ;
        RECT 4.000 2553.720 3515.600 2555.120 ;
        RECT 4.000 2508.200 3516.000 2553.720 ;
        RECT 4.400 2506.800 3516.000 2508.200 ;
        RECT 4.000 2485.760 3516.000 2506.800 ;
        RECT 4.000 2484.360 3515.600 2485.760 ;
        RECT 4.000 2439.520 3516.000 2484.360 ;
        RECT 4.400 2438.120 3516.000 2439.520 ;
        RECT 4.000 2415.720 3516.000 2438.120 ;
        RECT 4.000 2414.320 3515.600 2415.720 ;
        RECT 4.000 2370.840 3516.000 2414.320 ;
        RECT 4.400 2369.440 3516.000 2370.840 ;
        RECT 4.000 2345.680 3516.000 2369.440 ;
        RECT 4.000 2344.280 3515.600 2345.680 ;
        RECT 4.000 2302.160 3516.000 2344.280 ;
        RECT 4.400 2300.760 3516.000 2302.160 ;
        RECT 4.000 2275.640 3516.000 2300.760 ;
        RECT 4.000 2274.240 3515.600 2275.640 ;
        RECT 4.000 2233.480 3516.000 2274.240 ;
        RECT 4.400 2232.080 3516.000 2233.480 ;
        RECT 4.000 2205.600 3516.000 2232.080 ;
        RECT 4.000 2204.200 3515.600 2205.600 ;
        RECT 4.000 2164.800 3516.000 2204.200 ;
        RECT 4.400 2163.400 3516.000 2164.800 ;
        RECT 4.000 2135.560 3516.000 2163.400 ;
        RECT 4.000 2134.160 3515.600 2135.560 ;
        RECT 4.000 2096.120 3516.000 2134.160 ;
        RECT 4.400 2094.720 3516.000 2096.120 ;
        RECT 4.000 2065.520 3516.000 2094.720 ;
        RECT 4.000 2064.120 3515.600 2065.520 ;
        RECT 4.000 2027.440 3516.000 2064.120 ;
        RECT 4.400 2026.040 3516.000 2027.440 ;
        RECT 4.000 1995.480 3516.000 2026.040 ;
        RECT 4.000 1994.080 3515.600 1995.480 ;
        RECT 4.000 1958.760 3516.000 1994.080 ;
        RECT 4.400 1957.360 3516.000 1958.760 ;
        RECT 4.000 1925.440 3516.000 1957.360 ;
        RECT 4.000 1924.040 3515.600 1925.440 ;
        RECT 4.000 1890.080 3516.000 1924.040 ;
        RECT 4.400 1888.680 3516.000 1890.080 ;
        RECT 4.000 1855.400 3516.000 1888.680 ;
        RECT 4.000 1854.000 3515.600 1855.400 ;
        RECT 4.000 1820.720 3516.000 1854.000 ;
        RECT 4.400 1819.320 3516.000 1820.720 ;
        RECT 4.000 1785.360 3516.000 1819.320 ;
        RECT 4.000 1783.960 3515.600 1785.360 ;
        RECT 4.000 1752.040 3516.000 1783.960 ;
        RECT 4.400 1750.640 3516.000 1752.040 ;
        RECT 4.000 1715.320 3516.000 1750.640 ;
        RECT 4.000 1713.920 3515.600 1715.320 ;
        RECT 4.000 1683.360 3516.000 1713.920 ;
        RECT 4.400 1681.960 3516.000 1683.360 ;
        RECT 4.000 1645.280 3516.000 1681.960 ;
        RECT 4.000 1643.880 3515.600 1645.280 ;
        RECT 4.000 1614.680 3516.000 1643.880 ;
        RECT 4.400 1613.280 3516.000 1614.680 ;
        RECT 4.000 1575.240 3516.000 1613.280 ;
        RECT 4.000 1573.840 3515.600 1575.240 ;
        RECT 4.000 1546.000 3516.000 1573.840 ;
        RECT 4.400 1544.600 3516.000 1546.000 ;
        RECT 4.000 1505.200 3516.000 1544.600 ;
        RECT 4.000 1503.800 3515.600 1505.200 ;
        RECT 4.000 1477.320 3516.000 1503.800 ;
        RECT 4.400 1475.920 3516.000 1477.320 ;
        RECT 4.000 1435.160 3516.000 1475.920 ;
        RECT 4.000 1433.760 3515.600 1435.160 ;
        RECT 4.000 1408.640 3516.000 1433.760 ;
        RECT 4.400 1407.240 3516.000 1408.640 ;
        RECT 4.000 1365.120 3516.000 1407.240 ;
        RECT 4.000 1363.720 3515.600 1365.120 ;
        RECT 4.000 1339.960 3516.000 1363.720 ;
        RECT 4.400 1338.560 3516.000 1339.960 ;
        RECT 4.000 1295.080 3516.000 1338.560 ;
        RECT 4.000 1293.680 3515.600 1295.080 ;
        RECT 4.000 1271.280 3516.000 1293.680 ;
        RECT 4.400 1269.880 3516.000 1271.280 ;
        RECT 4.000 1225.720 3516.000 1269.880 ;
        RECT 4.000 1224.320 3515.600 1225.720 ;
        RECT 4.000 1202.600 3516.000 1224.320 ;
        RECT 4.400 1201.200 3516.000 1202.600 ;
        RECT 4.000 1155.680 3516.000 1201.200 ;
        RECT 4.000 1154.280 3515.600 1155.680 ;
        RECT 4.000 1133.920 3516.000 1154.280 ;
        RECT 4.400 1132.520 3516.000 1133.920 ;
        RECT 4.000 1085.640 3516.000 1132.520 ;
        RECT 4.000 1084.240 3515.600 1085.640 ;
        RECT 4.000 1065.240 3516.000 1084.240 ;
        RECT 4.400 1063.840 3516.000 1065.240 ;
        RECT 4.000 1015.600 3516.000 1063.840 ;
        RECT 4.000 1014.200 3515.600 1015.600 ;
        RECT 4.000 996.560 3516.000 1014.200 ;
        RECT 4.400 995.160 3516.000 996.560 ;
        RECT 4.000 945.560 3516.000 995.160 ;
        RECT 4.000 944.160 3515.600 945.560 ;
        RECT 4.000 927.880 3516.000 944.160 ;
        RECT 4.400 926.480 3516.000 927.880 ;
        RECT 4.000 875.520 3516.000 926.480 ;
        RECT 4.000 874.120 3515.600 875.520 ;
        RECT 4.000 859.200 3516.000 874.120 ;
        RECT 4.400 857.800 3516.000 859.200 ;
        RECT 4.000 805.480 3516.000 857.800 ;
        RECT 4.000 804.080 3515.600 805.480 ;
        RECT 4.000 790.520 3516.000 804.080 ;
        RECT 4.400 789.120 3516.000 790.520 ;
        RECT 4.000 735.440 3516.000 789.120 ;
        RECT 4.000 734.040 3515.600 735.440 ;
        RECT 4.000 721.840 3516.000 734.040 ;
        RECT 4.400 720.440 3516.000 721.840 ;
        RECT 4.000 665.400 3516.000 720.440 ;
        RECT 4.000 664.000 3515.600 665.400 ;
        RECT 4.000 653.160 3516.000 664.000 ;
        RECT 4.400 651.760 3516.000 653.160 ;
        RECT 4.000 595.360 3516.000 651.760 ;
        RECT 4.000 593.960 3515.600 595.360 ;
        RECT 4.000 584.480 3516.000 593.960 ;
        RECT 4.400 583.080 3516.000 584.480 ;
        RECT 4.000 525.320 3516.000 583.080 ;
        RECT 4.000 523.920 3515.600 525.320 ;
        RECT 4.000 515.800 3516.000 523.920 ;
        RECT 4.400 514.400 3516.000 515.800 ;
        RECT 4.000 455.280 3516.000 514.400 ;
        RECT 4.000 453.880 3515.600 455.280 ;
        RECT 4.000 447.120 3516.000 453.880 ;
        RECT 4.400 445.720 3516.000 447.120 ;
        RECT 4.000 385.240 3516.000 445.720 ;
        RECT 4.000 383.840 3515.600 385.240 ;
        RECT 4.000 378.440 3516.000 383.840 ;
        RECT 4.400 377.040 3516.000 378.440 ;
        RECT 4.000 315.200 3516.000 377.040 ;
        RECT 4.000 313.800 3515.600 315.200 ;
        RECT 4.000 309.760 3516.000 313.800 ;
        RECT 4.400 308.360 3516.000 309.760 ;
        RECT 4.000 245.160 3516.000 308.360 ;
        RECT 4.000 243.760 3515.600 245.160 ;
        RECT 4.000 241.080 3516.000 243.760 ;
        RECT 4.400 239.680 3516.000 241.080 ;
        RECT 4.000 175.120 3516.000 239.680 ;
        RECT 4.000 173.720 3515.600 175.120 ;
        RECT 4.000 172.400 3516.000 173.720 ;
        RECT 4.400 171.000 3516.000 172.400 ;
        RECT 4.000 105.080 3516.000 171.000 ;
        RECT 4.000 103.720 3515.600 105.080 ;
        RECT 4.400 103.680 3515.600 103.720 ;
        RECT 4.400 102.320 3516.000 103.680 ;
        RECT 4.000 35.720 3516.000 102.320 ;
        RECT 4.000 35.040 3515.600 35.720 ;
        RECT 4.400 34.320 3515.600 35.040 ;
        RECT 4.400 33.640 3516.000 34.320 ;
        RECT 4.000 16.495 3516.000 33.640 ;
      LAYER met4 ;
        RECT 350.000 440.000 3170.260 3659.800 ;
      LAYER met5 ;
        RECT -42.880 3744.880 -39.880 3744.890 ;
        RECT 3559.800 3744.880 3562.800 3744.890 ;
        RECT -42.880 3741.870 -39.880 3741.880 ;
        RECT 3559.800 3741.870 3562.800 3741.880 ;
        RECT -38.180 3740.180 -35.180 3740.190 ;
        RECT 3555.100 3740.180 3558.100 3740.190 ;
        RECT -38.180 3737.170 -35.180 3737.180 ;
        RECT 3555.100 3737.170 3558.100 3737.180 ;
        RECT -33.480 3735.480 -30.480 3735.490 ;
        RECT 3550.400 3735.480 3553.400 3735.490 ;
        RECT -33.480 3732.470 -30.480 3732.480 ;
        RECT 3550.400 3732.470 3553.400 3732.480 ;
        RECT -28.780 3730.780 -25.780 3730.790 ;
        RECT 3545.700 3730.780 3548.700 3730.790 ;
        RECT -28.780 3727.770 -25.780 3727.780 ;
        RECT 3545.700 3727.770 3548.700 3727.780 ;
        RECT -24.080 3726.080 -21.080 3726.090 ;
        RECT 3541.000 3726.080 3544.000 3726.090 ;
        RECT -24.080 3723.070 -21.080 3723.080 ;
        RECT 3541.000 3723.070 3544.000 3723.080 ;
        RECT -19.380 3721.380 -16.380 3721.390 ;
        RECT 3536.300 3721.380 3539.300 3721.390 ;
        RECT -19.380 3718.370 -16.380 3718.380 ;
        RECT 3536.300 3718.370 3539.300 3718.380 ;
        RECT -14.680 3716.680 -11.680 3716.690 ;
        RECT 94.020 3716.680 97.020 3716.690 ;
        RECT 274.020 3716.680 277.020 3716.690 ;
        RECT 454.020 3716.680 457.020 3716.690 ;
        RECT 634.020 3716.680 637.020 3716.690 ;
        RECT 814.020 3716.680 817.020 3716.690 ;
        RECT 994.020 3716.680 997.020 3716.690 ;
        RECT 1174.020 3716.680 1177.020 3716.690 ;
        RECT 1354.020 3716.680 1357.020 3716.690 ;
        RECT 1534.020 3716.680 1537.020 3716.690 ;
        RECT 1714.020 3716.680 1717.020 3716.690 ;
        RECT 1894.020 3716.680 1897.020 3716.690 ;
        RECT 2074.020 3716.680 2077.020 3716.690 ;
        RECT 2254.020 3716.680 2257.020 3716.690 ;
        RECT 2434.020 3716.680 2437.020 3716.690 ;
        RECT 2614.020 3716.680 2617.020 3716.690 ;
        RECT 2794.020 3716.680 2797.020 3716.690 ;
        RECT 2974.020 3716.680 2977.020 3716.690 ;
        RECT 3154.020 3716.680 3157.020 3716.690 ;
        RECT 3334.020 3716.680 3337.020 3716.690 ;
        RECT 3531.600 3716.680 3534.600 3716.690 ;
        RECT -14.680 3713.670 -11.680 3713.680 ;
        RECT 94.020 3713.670 97.020 3713.680 ;
        RECT 274.020 3713.670 277.020 3713.680 ;
        RECT 454.020 3713.670 457.020 3713.680 ;
        RECT 634.020 3713.670 637.020 3713.680 ;
        RECT 814.020 3713.670 817.020 3713.680 ;
        RECT 994.020 3713.670 997.020 3713.680 ;
        RECT 1174.020 3713.670 1177.020 3713.680 ;
        RECT 1354.020 3713.670 1357.020 3713.680 ;
        RECT 1534.020 3713.670 1537.020 3713.680 ;
        RECT 1714.020 3713.670 1717.020 3713.680 ;
        RECT 1894.020 3713.670 1897.020 3713.680 ;
        RECT 2074.020 3713.670 2077.020 3713.680 ;
        RECT 2254.020 3713.670 2257.020 3713.680 ;
        RECT 2434.020 3713.670 2437.020 3713.680 ;
        RECT 2614.020 3713.670 2617.020 3713.680 ;
        RECT 2794.020 3713.670 2797.020 3713.680 ;
        RECT 2974.020 3713.670 2977.020 3713.680 ;
        RECT 3154.020 3713.670 3157.020 3713.680 ;
        RECT 3334.020 3713.670 3337.020 3713.680 ;
        RECT 3531.600 3713.670 3534.600 3713.680 ;
        RECT -9.980 3711.980 -6.980 3711.990 ;
        RECT 4.020 3711.980 7.020 3711.990 ;
        RECT 184.020 3711.980 187.020 3711.990 ;
        RECT 364.020 3711.980 367.020 3711.990 ;
        RECT 544.020 3711.980 547.020 3711.990 ;
        RECT 724.020 3711.980 727.020 3711.990 ;
        RECT 904.020 3711.980 907.020 3711.990 ;
        RECT 1084.020 3711.980 1087.020 3711.990 ;
        RECT 1264.020 3711.980 1267.020 3711.990 ;
        RECT 1444.020 3711.980 1447.020 3711.990 ;
        RECT 1624.020 3711.980 1627.020 3711.990 ;
        RECT 1804.020 3711.980 1807.020 3711.990 ;
        RECT 1984.020 3711.980 1987.020 3711.990 ;
        RECT 2164.020 3711.980 2167.020 3711.990 ;
        RECT 2344.020 3711.980 2347.020 3711.990 ;
        RECT 2524.020 3711.980 2527.020 3711.990 ;
        RECT 2704.020 3711.980 2707.020 3711.990 ;
        RECT 2884.020 3711.980 2887.020 3711.990 ;
        RECT 3064.020 3711.980 3067.020 3711.990 ;
        RECT 3244.020 3711.980 3247.020 3711.990 ;
        RECT 3424.020 3711.980 3427.020 3711.990 ;
        RECT 3526.900 3711.980 3529.900 3711.990 ;
        RECT -9.980 3708.970 -6.980 3708.980 ;
        RECT 3526.900 3708.970 3529.900 3708.980 ;
        RECT 0.000 3613.980 3520.000 3707.380 ;
        RECT -9.980 3612.380 -6.980 3612.390 ;
        RECT 3526.900 3612.380 3529.900 3612.390 ;
        RECT -9.980 3609.370 -6.980 3609.380 ;
        RECT 3526.900 3609.370 3529.900 3609.380 ;
        RECT 0.000 3523.980 3520.000 3607.780 ;
        RECT -14.680 3522.380 -11.680 3522.390 ;
        RECT 3531.600 3522.380 3534.600 3522.390 ;
        RECT -14.680 3519.370 -11.680 3519.380 ;
        RECT 3531.600 3519.370 3534.600 3519.380 ;
        RECT 0.000 3433.980 3520.000 3517.780 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 3526.900 3432.380 3529.900 3432.390 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 3526.900 3429.370 3529.900 3429.380 ;
        RECT 0.000 3343.980 3520.000 3427.780 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 3531.600 3342.380 3534.600 3342.390 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 3531.600 3339.370 3534.600 3339.380 ;
        RECT 0.000 3253.980 3520.000 3337.780 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 3526.900 3252.380 3529.900 3252.390 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 3526.900 3249.370 3529.900 3249.380 ;
        RECT 0.000 3163.980 3520.000 3247.780 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 3531.600 3162.380 3534.600 3162.390 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 3531.600 3159.370 3534.600 3159.380 ;
        RECT 0.000 3073.980 3520.000 3157.780 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 3526.900 3072.380 3529.900 3072.390 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 3526.900 3069.370 3529.900 3069.380 ;
        RECT 0.000 2983.980 3520.000 3067.780 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 3531.600 2982.380 3534.600 2982.390 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 3531.600 2979.370 3534.600 2979.380 ;
        RECT 0.000 2893.980 3520.000 2977.780 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 3526.900 2892.380 3529.900 2892.390 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 3526.900 2889.370 3529.900 2889.380 ;
        RECT 0.000 2803.980 3520.000 2887.780 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 3531.600 2802.380 3534.600 2802.390 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 3531.600 2799.370 3534.600 2799.380 ;
        RECT 0.000 2713.980 3520.000 2797.780 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 3526.900 2712.380 3529.900 2712.390 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 3526.900 2709.370 3529.900 2709.380 ;
        RECT 0.000 2623.980 3520.000 2707.780 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 3531.600 2622.380 3534.600 2622.390 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 3531.600 2619.370 3534.600 2619.380 ;
        RECT 0.000 2533.980 3520.000 2617.780 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 3526.900 2532.380 3529.900 2532.390 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 3526.900 2529.370 3529.900 2529.380 ;
        RECT 0.000 2443.980 3520.000 2527.780 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 3531.600 2442.380 3534.600 2442.390 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 3531.600 2439.370 3534.600 2439.380 ;
        RECT 0.000 2353.980 3520.000 2437.780 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 3526.900 2352.380 3529.900 2352.390 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 3526.900 2349.370 3529.900 2349.380 ;
        RECT 0.000 2263.980 3520.000 2347.780 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 3531.600 2262.380 3534.600 2262.390 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 3531.600 2259.370 3534.600 2259.380 ;
        RECT 0.000 2173.980 3520.000 2257.780 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 3526.900 2172.380 3529.900 2172.390 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 3526.900 2169.370 3529.900 2169.380 ;
        RECT 0.000 2083.980 3520.000 2167.780 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 3531.600 2082.380 3534.600 2082.390 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 3531.600 2079.370 3534.600 2079.380 ;
        RECT 0.000 1993.980 3520.000 2077.780 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 3526.900 1992.380 3529.900 1992.390 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 3526.900 1989.370 3529.900 1989.380 ;
        RECT 0.000 1903.980 3520.000 1987.780 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 3531.600 1902.380 3534.600 1902.390 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 3531.600 1899.370 3534.600 1899.380 ;
        RECT 0.000 1813.980 3520.000 1897.780 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 3526.900 1812.380 3529.900 1812.390 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 3526.900 1809.370 3529.900 1809.380 ;
        RECT 0.000 1723.980 3520.000 1807.780 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 3531.600 1722.380 3534.600 1722.390 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 3531.600 1719.370 3534.600 1719.380 ;
        RECT 0.000 1633.980 3520.000 1717.780 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 3526.900 1632.380 3529.900 1632.390 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 3526.900 1629.370 3529.900 1629.380 ;
        RECT 0.000 1543.980 3520.000 1627.780 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 3531.600 1542.380 3534.600 1542.390 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 3531.600 1539.370 3534.600 1539.380 ;
        RECT 0.000 1453.980 3520.000 1537.780 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 3526.900 1452.380 3529.900 1452.390 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 3526.900 1449.370 3529.900 1449.380 ;
        RECT 0.000 1363.980 3520.000 1447.780 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 3531.600 1362.380 3534.600 1362.390 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 3531.600 1359.370 3534.600 1359.380 ;
        RECT 0.000 1273.980 3520.000 1357.780 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 3526.900 1272.380 3529.900 1272.390 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 3526.900 1269.370 3529.900 1269.380 ;
        RECT 0.000 1183.980 3520.000 1267.780 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 3531.600 1182.380 3534.600 1182.390 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 3531.600 1179.370 3534.600 1179.380 ;
        RECT 0.000 1093.980 3520.000 1177.780 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 3526.900 1092.380 3529.900 1092.390 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 3526.900 1089.370 3529.900 1089.380 ;
        RECT 0.000 1003.980 3520.000 1087.780 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 3531.600 1002.380 3534.600 1002.390 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 3531.600 999.370 3534.600 999.380 ;
        RECT 0.000 913.980 3520.000 997.780 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 3526.900 912.380 3529.900 912.390 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 3526.900 909.370 3529.900 909.380 ;
        RECT 0.000 823.980 3520.000 907.780 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 3531.600 822.380 3534.600 822.390 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 3531.600 819.370 3534.600 819.380 ;
        RECT 0.000 733.980 3520.000 817.780 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 3526.900 732.380 3529.900 732.390 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 3526.900 729.370 3529.900 729.380 ;
        RECT 0.000 643.980 3520.000 727.780 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 3531.600 642.380 3534.600 642.390 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 3531.600 639.370 3534.600 639.380 ;
        RECT 0.000 553.980 3520.000 637.780 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 3526.900 552.380 3529.900 552.390 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 3526.900 549.370 3529.900 549.380 ;
        RECT 0.000 463.980 3520.000 547.780 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 3531.600 462.380 3534.600 462.390 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 3531.600 459.370 3534.600 459.380 ;
        RECT 0.000 373.980 3520.000 457.780 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 3526.900 372.380 3529.900 372.390 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 3526.900 369.370 3529.900 369.380 ;
        RECT 0.000 283.980 3520.000 367.780 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 3531.600 282.380 3534.600 282.390 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 3531.600 279.370 3534.600 279.380 ;
        RECT 0.000 193.980 3520.000 277.780 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 3526.900 192.380 3529.900 192.390 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 3526.900 189.370 3529.900 189.380 ;
        RECT 0.000 103.980 3520.000 187.780 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 3531.600 102.380 3534.600 102.390 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 3531.600 99.370 3534.600 99.380 ;
        RECT 0.000 13.980 3520.000 97.780 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 3526.900 12.380 3529.900 12.390 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 3526.900 9.370 3529.900 9.380 ;
        RECT 0.000 0.000 3520.000 7.780 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 3064.020 -1.620 3067.020 -1.610 ;
        RECT 3244.020 -1.620 3247.020 -1.610 ;
        RECT 3424.020 -1.620 3427.020 -1.610 ;
        RECT 3526.900 -1.620 3529.900 -1.610 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 3064.020 -4.630 3067.020 -4.620 ;
        RECT 3244.020 -4.630 3247.020 -4.620 ;
        RECT 3424.020 -4.630 3427.020 -4.620 ;
        RECT 3526.900 -4.630 3529.900 -4.620 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2974.020 -6.320 2977.020 -6.310 ;
        RECT 3154.020 -6.320 3157.020 -6.310 ;
        RECT 3334.020 -6.320 3337.020 -6.310 ;
        RECT 3531.600 -6.320 3534.600 -6.310 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2974.020 -9.330 2977.020 -9.320 ;
        RECT 3154.020 -9.330 3157.020 -9.320 ;
        RECT 3334.020 -9.330 3337.020 -9.320 ;
        RECT 3531.600 -9.330 3534.600 -9.320 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 3536.300 -11.020 3539.300 -11.010 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 3536.300 -14.030 3539.300 -14.020 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 3541.000 -15.720 3544.000 -15.710 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 3541.000 -18.730 3544.000 -18.720 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 3545.700 -20.420 3548.700 -20.410 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 3545.700 -23.430 3548.700 -23.420 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 3550.400 -25.120 3553.400 -25.110 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 3550.400 -28.130 3553.400 -28.120 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 3555.100 -29.820 3558.100 -29.810 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 3555.100 -32.830 3558.100 -32.820 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 3559.800 -34.520 3562.800 -34.510 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 3559.800 -37.530 3562.800 -37.520 ;
  END
END user_project_wrapper
END LIBRARY

