##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Thu Dec 30 17:02:00 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 1120.100000 BY 919.700000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.200000 0.000000 2.340000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540000 0.000000 1.680000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.220000 0.000000 236.360000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.450000 0.000000 79.590000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.490000 0.000000 238.630000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.945000 0.000000 234.085000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.675000 0.000000 231.815000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.400000 0.000000 229.540000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.130000 0.000000 227.270000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.155000 0.000000 152.295000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.880000 0.000000 150.020000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.610000 0.000000 147.750000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.340000 0.000000 145.480000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.065000 0.000000 143.205000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.795000 0.000000 140.935000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.520000 0.000000 138.660000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250000 0.000000 136.390000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.980000 0.000000 134.120000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.705000 0.000000 131.845000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.435000 0.000000 129.575000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.160000 0.000000 127.300000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.890000 0.000000 125.030000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.620000 0.000000 122.760000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.345000 0.000000 120.485000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.075000 0.000000 118.215000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.800000 0.000000 115.940000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.530000 0.000000 113.670000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.260000 0.000000 111.400000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.985000 0.000000 109.125000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.715000 0.000000 106.855000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.440000 0.000000 104.580000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.170000 0.000000 102.310000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.900000 0.000000 100.040000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.625000 0.000000 97.765000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.355000 0.000000 95.495000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080000 0.000000 93.220000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.810000 0.000000 90.950000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.540000 0.000000 88.680000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.265000 0.000000 86.405000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.995000 0.000000 84.135000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.720000 0.000000 81.860000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.180000 0.000000 77.320000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.905000 0.000000 75.045000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.635000 0.000000 72.775000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.360000 0.000000 70.500000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.090000 0.000000 68.230000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.820000 0.000000 65.960000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.545000 0.000000 63.685000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.275000 0.000000 61.415000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.000000 0.000000 59.140000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.730000 0.000000 56.870000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.460000 0.000000 54.600000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.185000 0.000000 52.325000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.915000 0.000000 50.055000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.640000 0.000000 47.780000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.370000 0.000000 45.510000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.100000 0.000000 43.240000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.825000 0.000000 40.965000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.555000 0.000000 38.695000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.280000 0.000000 36.420000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.010000 0.000000 34.150000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.740000 0.000000 31.880000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.465000 0.000000 29.605000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.195000 0.000000 27.335000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.920000 0.000000 25.060000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.650000 0.000000 22.790000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.380000 0.000000 20.520000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.105000 0.000000 18.245000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.835000 0.000000 15.975000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.560000 0.000000 13.700000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.290000 0.000000 11.430000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.020000 0.000000 9.160000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.745000 0.000000 6.885000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.475000 0.000000 4.615000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.860000 0.000000 225.000000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.585000 0.000000 222.725000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.315000 0.000000 220.455000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.040000 0.000000 218.180000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.770000 0.000000 215.910000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.500000 0.000000 213.640000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.225000 0.000000 211.365000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.955000 0.000000 209.095000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.680000 0.000000 206.820000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.410000 0.000000 204.550000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.140000 0.000000 202.280000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.865000 0.000000 200.005000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.595000 0.000000 197.735000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.320000 0.000000 195.460000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.050000 0.000000 193.190000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.780000 0.000000 190.920000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.505000 0.000000 188.645000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.235000 0.000000 186.375000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.960000 0.000000 184.100000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.690000 0.000000 181.830000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.420000 0.000000 179.560000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.145000 0.000000 177.285000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.875000 0.000000 175.015000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.600000 0.000000 172.740000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.330000 0.000000 170.470000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060000 0.000000 168.200000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.785000 0.000000 165.925000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.515000 0.000000 163.655000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.240000 0.000000 161.380000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.970000 0.000000 159.110000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.700000 0.000000 156.840000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.425000 0.000000 154.565000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.305000 0.000000 529.445000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.035000 0.000000 527.175000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.760000 0.000000 524.900000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.490000 0.000000 522.630000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.220000 0.000000 520.360000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.945000 0.000000 518.085000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.675000 0.000000 515.815000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.400000 0.000000 513.540000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.130000 0.000000 511.270000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.860000 0.000000 509.000000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.585000 0.000000 506.725000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.315000 0.000000 504.455000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.040000 0.000000 502.180000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.770000 0.000000 499.910000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.500000 0.000000 497.640000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.225000 0.000000 495.365000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.955000 0.000000 493.095000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.680000 0.000000 490.820000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.410000 0.000000 488.550000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.140000 0.000000 486.280000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.865000 0.000000 484.005000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.595000 0.000000 481.735000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.320000 0.000000 479.460000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.050000 0.000000 477.190000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.780000 0.000000 474.920000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.505000 0.000000 472.645000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.235000 0.000000 470.375000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.960000 0.000000 468.100000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.690000 0.000000 465.830000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.420000 0.000000 463.560000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.145000 0.000000 461.285000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.875000 0.000000 459.015000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.600000 0.000000 456.740000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.330000 0.000000 454.470000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.060000 0.000000 452.200000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.785000 0.000000 449.925000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.515000 0.000000 447.655000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.240000 0.000000 445.380000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.970000 0.000000 443.110000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.700000 0.000000 440.840000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.425000 0.000000 438.565000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.155000 0.000000 436.295000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.880000 0.000000 434.020000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.610000 0.000000 431.750000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.340000 0.000000 429.480000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.065000 0.000000 427.205000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.795000 0.000000 424.935000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.520000 0.000000 422.660000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.250000 0.000000 420.390000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.980000 0.000000 418.120000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.705000 0.000000 415.845000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.435000 0.000000 413.575000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.160000 0.000000 411.300000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.890000 0.000000 409.030000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.620000 0.000000 406.760000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.345000 0.000000 404.485000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.075000 0.000000 402.215000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.800000 0.000000 399.940000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530000 0.000000 397.670000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.260000 0.000000 395.400000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.985000 0.000000 393.125000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.715000 0.000000 390.855000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.440000 0.000000 388.580000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.170000 0.000000 386.310000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.900000 0.000000 384.040000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.625000 0.000000 381.765000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.355000 0.000000 379.495000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.080000 0.000000 377.220000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.810000 0.000000 374.950000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.540000 0.000000 372.680000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.265000 0.000000 370.405000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.995000 0.000000 368.135000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.720000 0.000000 365.860000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.450000 0.000000 363.590000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.180000 0.000000 361.320000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.905000 0.000000 359.045000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.635000 0.000000 356.775000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.360000 0.000000 354.500000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.090000 0.000000 352.230000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.820000 0.000000 349.960000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.545000 0.000000 347.685000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.275000 0.000000 345.415000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.000000 0.000000 343.140000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.730000 0.000000 340.870000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.460000 0.000000 338.600000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.185000 0.000000 336.325000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.915000 0.000000 334.055000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.640000 0.000000 331.780000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.370000 0.000000 329.510000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.100000 0.000000 327.240000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.825000 0.000000 324.965000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.555000 0.000000 322.695000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.280000 0.000000 320.420000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.010000 0.000000 318.150000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.740000 0.000000 315.880000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.465000 0.000000 313.605000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.195000 0.000000 311.335000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.920000 0.000000 309.060000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.650000 0.000000 306.790000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.380000 0.000000 304.520000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.105000 0.000000 302.245000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.835000 0.000000 299.975000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.560000 0.000000 297.700000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.290000 0.000000 295.430000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.020000 0.000000 293.160000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.745000 0.000000 290.885000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.475000 0.000000 288.615000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.200000 0.000000 286.340000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.930000 0.000000 284.070000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.660000 0.000000 281.800000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.385000 0.000000 279.525000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.115000 0.000000 277.255000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.840000 0.000000 274.980000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.570000 0.000000 272.710000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.300000 0.000000 270.440000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.025000 0.000000 268.165000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.755000 0.000000 265.895000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.480000 0.000000 263.620000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.210000 0.000000 261.350000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.940000 0.000000 259.080000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.665000 0.000000 256.805000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.395000 0.000000 254.535000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.120000 0.000000 252.260000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.850000 0.000000 249.990000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.580000 0.000000 247.720000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.305000 0.000000 245.445000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.035000 0.000000 243.175000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.760000 0.000000 240.900000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.120000 0.000000 820.260000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.850000 0.000000 817.990000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.580000 0.000000 815.720000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.305000 0.000000 813.445000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.035000 0.000000 811.175000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.760000 0.000000 808.900000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.490000 0.000000 806.630000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.220000 0.000000 804.360000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.945000 0.000000 802.085000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.675000 0.000000 799.815000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.400000 0.000000 797.540000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.130000 0.000000 795.270000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.860000 0.000000 793.000000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.585000 0.000000 790.725000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.315000 0.000000 788.455000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.040000 0.000000 786.180000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.770000 0.000000 783.910000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.500000 0.000000 781.640000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.225000 0.000000 779.365000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.955000 0.000000 777.095000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.680000 0.000000 774.820000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.410000 0.000000 772.550000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.140000 0.000000 770.280000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.865000 0.000000 768.005000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.595000 0.000000 765.735000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.320000 0.000000 763.460000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.050000 0.000000 761.190000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.780000 0.000000 758.920000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.505000 0.000000 756.645000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.235000 0.000000 754.375000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.960000 0.000000 752.100000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.690000 0.000000 749.830000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.420000 0.000000 747.560000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.145000 0.000000 745.285000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.875000 0.000000 743.015000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.600000 0.000000 740.740000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.330000 0.000000 738.470000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.060000 0.000000 736.200000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.785000 0.000000 733.925000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.515000 0.000000 731.655000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.240000 0.000000 729.380000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.970000 0.000000 727.110000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.700000 0.000000 724.840000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.425000 0.000000 722.565000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.155000 0.000000 720.295000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.880000 0.000000 718.020000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.610000 0.000000 715.750000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.340000 0.000000 713.480000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.065000 0.000000 711.205000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.795000 0.000000 708.935000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.520000 0.000000 706.660000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.250000 0.000000 704.390000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.980000 0.000000 702.120000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.705000 0.000000 699.845000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.435000 0.000000 697.575000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.160000 0.000000 695.300000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.890000 0.000000 693.030000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.620000 0.000000 690.760000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.345000 0.000000 688.485000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.075000 0.000000 686.215000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.800000 0.000000 683.940000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.530000 0.000000 681.670000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.260000 0.000000 679.400000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.985000 0.000000 677.125000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.715000 0.000000 674.855000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.440000 0.000000 672.580000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.170000 0.000000 670.310000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.900000 0.000000 668.040000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.625000 0.000000 665.765000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.355000 0.000000 663.495000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.080000 0.000000 661.220000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810000 0.000000 658.950000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.540000 0.000000 656.680000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.265000 0.000000 654.405000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.995000 0.000000 652.135000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.720000 0.000000 649.860000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.450000 0.000000 647.590000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.180000 0.000000 645.320000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.905000 0.000000 643.045000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.635000 0.000000 640.775000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.360000 0.000000 638.500000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.090000 0.000000 636.230000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.820000 0.000000 633.960000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.545000 0.000000 631.685000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.275000 0.000000 629.415000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.000000 0.000000 627.140000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.730000 0.000000 624.870000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.460000 0.000000 622.600000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.185000 0.000000 620.325000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.915000 0.000000 618.055000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.640000 0.000000 615.780000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.370000 0.000000 613.510000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.100000 0.000000 611.240000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.825000 0.000000 608.965000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.555000 0.000000 606.695000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.280000 0.000000 604.420000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.010000 0.000000 602.150000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.740000 0.000000 599.880000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.465000 0.000000 597.605000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.195000 0.000000 595.335000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.920000 0.000000 593.060000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.650000 0.000000 590.790000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.380000 0.000000 588.520000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.105000 0.000000 586.245000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.835000 0.000000 583.975000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.560000 0.000000 581.700000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.290000 0.000000 579.430000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.020000 0.000000 577.160000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.745000 0.000000 574.885000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.475000 0.000000 572.615000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.200000 0.000000 570.340000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.930000 0.000000 568.070000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.660000 0.000000 565.800000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.385000 0.000000 563.525000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.115000 0.000000 561.255000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.840000 0.000000 558.980000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.570000 0.000000 556.710000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.300000 0.000000 554.440000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.025000 0.000000 552.165000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.755000 0.000000 549.895000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.480000 0.000000 547.620000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.210000 0.000000 545.350000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.940000 0.000000 543.080000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.665000 0.000000 540.805000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.395000 0.000000 538.535000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.120000 0.000000 536.260000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.850000 0.000000 533.990000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.580000 0.000000 531.720000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.940000 0.000000 1111.080000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.665000 0.000000 1108.805000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.395000 0.000000 1106.535000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.120000 0.000000 1104.260000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.850000 0.000000 1101.990000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.580000 0.000000 1099.720000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.305000 0.000000 1097.445000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.035000 0.000000 1095.175000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.760000 0.000000 1092.900000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.490000 0.000000 1090.630000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.220000 0.000000 1088.360000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.945000 0.000000 1086.085000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.675000 0.000000 1083.815000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.400000 0.000000 1081.540000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.130000 0.000000 1079.270000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.860000 0.000000 1077.000000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.585000 0.000000 1074.725000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.315000 0.000000 1072.455000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.040000 0.000000 1070.180000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.770000 0.000000 1067.910000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.500000 0.000000 1065.640000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.225000 0.000000 1063.365000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.955000 0.000000 1061.095000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.680000 0.000000 1058.820000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.410000 0.000000 1056.550000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.140000 0.000000 1054.280000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.865000 0.000000 1052.005000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.595000 0.000000 1049.735000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.320000 0.000000 1047.460000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.050000 0.000000 1045.190000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.780000 0.000000 1042.920000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.505000 0.000000 1040.645000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.235000 0.000000 1038.375000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.960000 0.000000 1036.100000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.690000 0.000000 1033.830000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.420000 0.000000 1031.560000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.145000 0.000000 1029.285000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.875000 0.000000 1027.015000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.600000 0.000000 1024.740000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.330000 0.000000 1022.470000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.060000 0.000000 1020.200000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.785000 0.000000 1017.925000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.515000 0.000000 1015.655000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.240000 0.000000 1013.380000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.970000 0.000000 1011.110000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.700000 0.000000 1008.840000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.425000 0.000000 1006.565000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.155000 0.000000 1004.295000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.880000 0.000000 1002.020000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.610000 0.000000 999.750000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.340000 0.000000 997.480000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.065000 0.000000 995.205000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.795000 0.000000 992.935000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.520000 0.000000 990.660000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.250000 0.000000 988.390000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.980000 0.000000 986.120000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.705000 0.000000 983.845000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.435000 0.000000 981.575000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.160000 0.000000 979.300000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.890000 0.000000 977.030000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.620000 0.000000 974.760000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.345000 0.000000 972.485000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.075000 0.000000 970.215000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.800000 0.000000 967.940000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.530000 0.000000 965.670000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.260000 0.000000 963.400000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.985000 0.000000 961.125000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.715000 0.000000 958.855000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.440000 0.000000 956.580000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.170000 0.000000 954.310000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.900000 0.000000 952.040000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.625000 0.000000 949.765000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.355000 0.000000 947.495000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.080000 0.000000 945.220000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.810000 0.000000 942.950000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.540000 0.000000 940.680000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.265000 0.000000 938.405000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.995000 0.000000 936.135000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.720000 0.000000 933.860000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.450000 0.000000 931.590000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.180000 0.000000 929.320000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.905000 0.000000 927.045000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.635000 0.000000 924.775000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.360000 0.000000 922.500000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090000 0.000000 920.230000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.820000 0.000000 917.960000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.545000 0.000000 915.685000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.275000 0.000000 913.415000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.000000 0.000000 911.140000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.730000 0.000000 908.870000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.460000 0.000000 906.600000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.185000 0.000000 904.325000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.915000 0.000000 902.055000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.640000 0.000000 899.780000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.370000 0.000000 897.510000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.100000 0.000000 895.240000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.825000 0.000000 892.965000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.555000 0.000000 890.695000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.280000 0.000000 888.420000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.010000 0.000000 886.150000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.740000 0.000000 883.880000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.465000 0.000000 881.605000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.195000 0.000000 879.335000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.920000 0.000000 877.060000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.650000 0.000000 874.790000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.380000 0.000000 872.520000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.105000 0.000000 870.245000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.835000 0.000000 867.975000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.560000 0.000000 865.700000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.290000 0.000000 863.430000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.020000 0.000000 861.160000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.745000 0.000000 858.885000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.475000 0.000000 856.615000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.200000 0.000000 854.340000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.930000 0.000000 852.070000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.660000 0.000000 849.800000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.385000 0.000000 847.525000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.115000 0.000000 845.255000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.840000 0.000000 842.980000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.570000 0.000000 840.710000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.300000 0.000000 838.440000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.025000 0.000000 836.165000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.755000 0.000000 833.895000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.480000 0.000000 831.620000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.210000 0.000000 829.350000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.940000 0.000000 827.080000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.665000 0.000000 824.805000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.395000 0.000000 822.535000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.555000 0.800000 34.855000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.610000 0.800000 86.910000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.665000 0.800000 138.965000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 208.075000 0.800000 208.375000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 277.480000 0.800000 277.780000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 346.890000 0.800000 347.190000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 416.300000 0.800000 416.600000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 485.705000 0.800000 486.005000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 555.115000 0.800000 555.415000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 624.520000 0.800000 624.820000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 693.930000 0.800000 694.230000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 763.340000 0.800000 763.640000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 832.745000 0.800000 833.045000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 902.155000 0.800000 902.455000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.935000 919.210000 96.075000 919.700000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.945000 919.210000 224.085000 919.700000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.950000 919.210000 352.090000 919.700000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.960000 919.210000 480.100000 919.700000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.970000 919.210000 608.110000 919.700000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.975000 919.210000 736.115000 919.700000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.985000 919.210000 864.125000 919.700000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.990000 919.210000 992.130000 919.700000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.960000 919.210000 1118.100000 919.700000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 884.150000 1120.100000 884.450000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 813.405000 1120.100000 813.705000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 742.660000 1120.100000 742.960000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 671.920000 1120.100000 672.220000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 601.175000 1120.100000 601.475000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 530.430000 1120.100000 530.730000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 459.685000 1120.100000 459.985000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 388.940000 1120.100000 389.240000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 318.200000 1120.100000 318.500000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 265.140000 1120.100000 265.440000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 212.080000 1120.100000 212.380000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 159.025000 1120.100000 159.325000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 105.965000 1120.100000 106.265000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 52.910000 1120.100000 53.210000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 2.560000 1120.100000 2.860000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.200000 0.800000 17.500000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 69.260000 0.800000 69.560000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 121.315000 0.800000 121.615000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 190.720000 0.800000 191.020000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 260.130000 0.800000 260.430000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 329.540000 0.800000 329.840000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 398.945000 0.800000 399.245000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 468.355000 0.800000 468.655000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 537.760000 0.800000 538.060000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 607.170000 0.800000 607.470000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 676.580000 0.800000 676.880000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 745.985000 0.800000 746.285000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 815.395000 0.800000 815.695000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 884.800000 0.800000 885.100000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.935000 919.210000 64.075000 919.700000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.940000 919.210000 192.080000 919.700000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.950000 919.210000 320.090000 919.700000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.960000 919.210000 448.100000 919.700000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.965000 919.210000 576.105000 919.700000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.975000 919.210000 704.115000 919.700000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.980000 919.210000 832.120000 919.700000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.990000 919.210000 960.130000 919.700000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.000000 919.210000 1088.140000 919.700000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 901.835000 1120.100000 902.135000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 831.090000 1120.100000 831.390000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 760.350000 1120.100000 760.650000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 689.605000 1120.100000 689.905000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 618.860000 1120.100000 619.160000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 548.115000 1120.100000 548.415000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 477.370000 1120.100000 477.670000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 406.630000 1120.100000 406.930000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 335.885000 1120.100000 336.185000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 282.825000 1120.100000 283.125000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 229.770000 1120.100000 230.070000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 176.710000 1120.100000 177.010000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 123.650000 1120.100000 123.950000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 70.595000 1120.100000 70.895000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 17.535000 1120.100000 17.835000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 3.170000 0.800000 3.470000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 51.905000 0.800000 52.205000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.960000 0.800000 104.260000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 173.370000 0.800000 173.670000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 242.780000 0.800000 243.080000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 312.185000 0.800000 312.485000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 381.595000 0.800000 381.895000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 451.000000 0.800000 451.300000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 520.410000 0.800000 520.710000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 589.820000 0.800000 590.120000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 659.225000 0.800000 659.525000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 728.635000 0.800000 728.935000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 798.040000 0.800000 798.340000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 867.450000 0.800000 867.750000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.930000 919.210000 32.070000 919.700000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.940000 919.210000 160.080000 919.700000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.950000 919.210000 288.090000 919.700000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.955000 919.210000 416.095000 919.700000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.965000 919.210000 544.105000 919.700000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.970000 919.210000 672.110000 919.700000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.980000 919.210000 800.120000 919.700000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.990000 919.210000 928.130000 919.700000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.995000 919.210000 1056.135000 919.700000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 915.730000 1120.100000 916.030000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 848.780000 1120.100000 849.080000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 778.035000 1120.100000 778.335000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 707.290000 1120.100000 707.590000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 636.545000 1120.100000 636.845000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 565.800000 1120.100000 566.100000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 495.060000 1120.100000 495.360000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 424.315000 1120.100000 424.615000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 353.570000 1120.100000 353.870000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 300.510000 1120.100000 300.810000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 247.455000 1120.100000 247.755000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 194.395000 1120.100000 194.695000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 141.340000 1120.100000 141.640000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 88.280000 1120.100000 88.580000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 35.220000 1120.100000 35.520000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.020000 0.800000 156.320000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 225.425000 0.800000 225.725000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.835000 0.800000 295.135000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 364.240000 0.800000 364.540000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 433.650000 0.800000 433.950000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 503.060000 0.800000 503.360000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 572.465000 0.800000 572.765000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 641.875000 0.800000 642.175000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 711.280000 0.800000 711.580000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 780.690000 0.800000 780.990000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 850.100000 0.800000 850.400000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 916.340000 0.800000 916.640000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.940000 919.210000 128.080000 919.700000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.945000 919.210000 256.085000 919.700000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.955000 919.210000 384.095000 919.700000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.960000 919.210000 512.100000 919.700000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.970000 919.210000 640.110000 919.700000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.980000 919.210000 768.120000 919.700000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.985000 919.210000 896.125000 919.700000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.995000 919.210000 1024.135000 919.700000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000000 919.210000 2.140000 919.700000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 866.465000 1120.100000 866.765000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 795.720000 1120.100000 796.020000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 724.975000 1120.100000 725.275000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 654.230000 1120.100000 654.530000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 583.490000 1120.100000 583.790000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 512.745000 1120.100000 513.045000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 442.000000 1120.100000 442.300000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.300000 371.255000 1120.100000 371.555000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.210000 0.000000 1113.350000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.580000 0.000000 1116.720000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.755000 0.000000 1117.895000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.480000 0.000000 1115.620000 0.490000 ;
    END
  END user_irq[0]
  PIN VWPR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.060000 1.930000 4.060000 916.580000 ;
    END
  END VWPR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1112.040000 5.930000 1114.040000 912.580000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 5.930000 8.060000 912.580000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 608.675000 493.280000 610.415000 888.060000 ;
      LAYER met4 ;
        RECT 1083.995000 493.280000 1085.735000 888.060000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 25.480000 489.805000 27.220000 884.585000 ;
      LAYER met4 ;
        RECT 500.800000 489.805000 502.540000 884.585000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1094.420000 27.325000 1096.160000 422.105000 ;
      LAYER met4 ;
        RECT 619.100000 27.325000 620.840000 422.105000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1116.040000 1.930000 1118.040000 916.580000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1080.595000 496.680000 1082.335000 884.660000 ;
      LAYER met4 ;
        RECT 612.075000 496.680000 613.815000 884.660000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 497.400000 493.205000 499.140000 881.185000 ;
      LAYER met4 ;
        RECT 28.880000 493.205000 30.620000 881.185000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 622.500000 30.725000 624.240000 418.705000 ;
      LAYER met4 ;
        RECT 1091.020000 30.725000 1092.760000 418.705000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1120.100000 919.700000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1120.100000 919.700000 ;
    LAYER met2 ;
      RECT 1118.240000 919.070000 1120.100000 919.700000 ;
      RECT 1088.280000 919.070000 1117.820000 919.700000 ;
      RECT 1056.275000 919.070000 1087.860000 919.700000 ;
      RECT 1024.275000 919.070000 1055.855000 919.700000 ;
      RECT 992.270000 919.070000 1023.855000 919.700000 ;
      RECT 960.270000 919.070000 991.850000 919.700000 ;
      RECT 928.270000 919.070000 959.850000 919.700000 ;
      RECT 896.265000 919.070000 927.850000 919.700000 ;
      RECT 864.265000 919.070000 895.845000 919.700000 ;
      RECT 832.260000 919.070000 863.845000 919.700000 ;
      RECT 800.260000 919.070000 831.840000 919.700000 ;
      RECT 768.260000 919.070000 799.840000 919.700000 ;
      RECT 736.255000 919.070000 767.840000 919.700000 ;
      RECT 704.255000 919.070000 735.835000 919.700000 ;
      RECT 672.250000 919.070000 703.835000 919.700000 ;
      RECT 640.250000 919.070000 671.830000 919.700000 ;
      RECT 608.250000 919.070000 639.830000 919.700000 ;
      RECT 576.245000 919.070000 607.830000 919.700000 ;
      RECT 544.245000 919.070000 575.825000 919.700000 ;
      RECT 512.240000 919.070000 543.825000 919.700000 ;
      RECT 480.240000 919.070000 511.820000 919.700000 ;
      RECT 448.240000 919.070000 479.820000 919.700000 ;
      RECT 416.235000 919.070000 447.820000 919.700000 ;
      RECT 384.235000 919.070000 415.815000 919.700000 ;
      RECT 352.230000 919.070000 383.815000 919.700000 ;
      RECT 320.230000 919.070000 351.810000 919.700000 ;
      RECT 288.230000 919.070000 319.810000 919.700000 ;
      RECT 256.225000 919.070000 287.810000 919.700000 ;
      RECT 224.225000 919.070000 255.805000 919.700000 ;
      RECT 192.220000 919.070000 223.805000 919.700000 ;
      RECT 160.220000 919.070000 191.800000 919.700000 ;
      RECT 128.220000 919.070000 159.800000 919.700000 ;
      RECT 96.215000 919.070000 127.800000 919.700000 ;
      RECT 64.215000 919.070000 95.795000 919.700000 ;
      RECT 32.210000 919.070000 63.795000 919.700000 ;
      RECT 2.280000 919.070000 31.790000 919.700000 ;
      RECT 0.000000 919.070000 1.860000 919.700000 ;
      RECT 0.000000 0.630000 1120.100000 919.070000 ;
      RECT 1118.035000 0.000000 1120.100000 0.630000 ;
      RECT 1116.860000 0.000000 1117.615000 0.630000 ;
      RECT 1115.760000 0.000000 1116.440000 0.630000 ;
      RECT 1113.490000 0.000000 1115.340000 0.630000 ;
      RECT 1111.220000 0.000000 1113.070000 0.630000 ;
      RECT 1108.945000 0.000000 1110.800000 0.630000 ;
      RECT 1106.675000 0.000000 1108.525000 0.630000 ;
      RECT 1104.400000 0.000000 1106.255000 0.630000 ;
      RECT 1102.130000 0.000000 1103.980000 0.630000 ;
      RECT 1099.860000 0.000000 1101.710000 0.630000 ;
      RECT 1097.585000 0.000000 1099.440000 0.630000 ;
      RECT 1095.315000 0.000000 1097.165000 0.630000 ;
      RECT 1093.040000 0.000000 1094.895000 0.630000 ;
      RECT 1090.770000 0.000000 1092.620000 0.630000 ;
      RECT 1088.500000 0.000000 1090.350000 0.630000 ;
      RECT 1086.225000 0.000000 1088.080000 0.630000 ;
      RECT 1083.955000 0.000000 1085.805000 0.630000 ;
      RECT 1081.680000 0.000000 1083.535000 0.630000 ;
      RECT 1079.410000 0.000000 1081.260000 0.630000 ;
      RECT 1077.140000 0.000000 1078.990000 0.630000 ;
      RECT 1074.865000 0.000000 1076.720000 0.630000 ;
      RECT 1072.595000 0.000000 1074.445000 0.630000 ;
      RECT 1070.320000 0.000000 1072.175000 0.630000 ;
      RECT 1068.050000 0.000000 1069.900000 0.630000 ;
      RECT 1065.780000 0.000000 1067.630000 0.630000 ;
      RECT 1063.505000 0.000000 1065.360000 0.630000 ;
      RECT 1061.235000 0.000000 1063.085000 0.630000 ;
      RECT 1058.960000 0.000000 1060.815000 0.630000 ;
      RECT 1056.690000 0.000000 1058.540000 0.630000 ;
      RECT 1054.420000 0.000000 1056.270000 0.630000 ;
      RECT 1052.145000 0.000000 1054.000000 0.630000 ;
      RECT 1049.875000 0.000000 1051.725000 0.630000 ;
      RECT 1047.600000 0.000000 1049.455000 0.630000 ;
      RECT 1045.330000 0.000000 1047.180000 0.630000 ;
      RECT 1043.060000 0.000000 1044.910000 0.630000 ;
      RECT 1040.785000 0.000000 1042.640000 0.630000 ;
      RECT 1038.515000 0.000000 1040.365000 0.630000 ;
      RECT 1036.240000 0.000000 1038.095000 0.630000 ;
      RECT 1033.970000 0.000000 1035.820000 0.630000 ;
      RECT 1031.700000 0.000000 1033.550000 0.630000 ;
      RECT 1029.425000 0.000000 1031.280000 0.630000 ;
      RECT 1027.155000 0.000000 1029.005000 0.630000 ;
      RECT 1024.880000 0.000000 1026.735000 0.630000 ;
      RECT 1022.610000 0.000000 1024.460000 0.630000 ;
      RECT 1020.340000 0.000000 1022.190000 0.630000 ;
      RECT 1018.065000 0.000000 1019.920000 0.630000 ;
      RECT 1015.795000 0.000000 1017.645000 0.630000 ;
      RECT 1013.520000 0.000000 1015.375000 0.630000 ;
      RECT 1011.250000 0.000000 1013.100000 0.630000 ;
      RECT 1008.980000 0.000000 1010.830000 0.630000 ;
      RECT 1006.705000 0.000000 1008.560000 0.630000 ;
      RECT 1004.435000 0.000000 1006.285000 0.630000 ;
      RECT 1002.160000 0.000000 1004.015000 0.630000 ;
      RECT 999.890000 0.000000 1001.740000 0.630000 ;
      RECT 997.620000 0.000000 999.470000 0.630000 ;
      RECT 995.345000 0.000000 997.200000 0.630000 ;
      RECT 993.075000 0.000000 994.925000 0.630000 ;
      RECT 990.800000 0.000000 992.655000 0.630000 ;
      RECT 988.530000 0.000000 990.380000 0.630000 ;
      RECT 986.260000 0.000000 988.110000 0.630000 ;
      RECT 983.985000 0.000000 985.840000 0.630000 ;
      RECT 981.715000 0.000000 983.565000 0.630000 ;
      RECT 979.440000 0.000000 981.295000 0.630000 ;
      RECT 977.170000 0.000000 979.020000 0.630000 ;
      RECT 974.900000 0.000000 976.750000 0.630000 ;
      RECT 972.625000 0.000000 974.480000 0.630000 ;
      RECT 970.355000 0.000000 972.205000 0.630000 ;
      RECT 968.080000 0.000000 969.935000 0.630000 ;
      RECT 965.810000 0.000000 967.660000 0.630000 ;
      RECT 963.540000 0.000000 965.390000 0.630000 ;
      RECT 961.265000 0.000000 963.120000 0.630000 ;
      RECT 958.995000 0.000000 960.845000 0.630000 ;
      RECT 956.720000 0.000000 958.575000 0.630000 ;
      RECT 954.450000 0.000000 956.300000 0.630000 ;
      RECT 952.180000 0.000000 954.030000 0.630000 ;
      RECT 949.905000 0.000000 951.760000 0.630000 ;
      RECT 947.635000 0.000000 949.485000 0.630000 ;
      RECT 945.360000 0.000000 947.215000 0.630000 ;
      RECT 943.090000 0.000000 944.940000 0.630000 ;
      RECT 940.820000 0.000000 942.670000 0.630000 ;
      RECT 938.545000 0.000000 940.400000 0.630000 ;
      RECT 936.275000 0.000000 938.125000 0.630000 ;
      RECT 934.000000 0.000000 935.855000 0.630000 ;
      RECT 931.730000 0.000000 933.580000 0.630000 ;
      RECT 929.460000 0.000000 931.310000 0.630000 ;
      RECT 927.185000 0.000000 929.040000 0.630000 ;
      RECT 924.915000 0.000000 926.765000 0.630000 ;
      RECT 922.640000 0.000000 924.495000 0.630000 ;
      RECT 920.370000 0.000000 922.220000 0.630000 ;
      RECT 918.100000 0.000000 919.950000 0.630000 ;
      RECT 915.825000 0.000000 917.680000 0.630000 ;
      RECT 913.555000 0.000000 915.405000 0.630000 ;
      RECT 911.280000 0.000000 913.135000 0.630000 ;
      RECT 909.010000 0.000000 910.860000 0.630000 ;
      RECT 906.740000 0.000000 908.590000 0.630000 ;
      RECT 904.465000 0.000000 906.320000 0.630000 ;
      RECT 902.195000 0.000000 904.045000 0.630000 ;
      RECT 899.920000 0.000000 901.775000 0.630000 ;
      RECT 897.650000 0.000000 899.500000 0.630000 ;
      RECT 895.380000 0.000000 897.230000 0.630000 ;
      RECT 893.105000 0.000000 894.960000 0.630000 ;
      RECT 890.835000 0.000000 892.685000 0.630000 ;
      RECT 888.560000 0.000000 890.415000 0.630000 ;
      RECT 886.290000 0.000000 888.140000 0.630000 ;
      RECT 884.020000 0.000000 885.870000 0.630000 ;
      RECT 881.745000 0.000000 883.600000 0.630000 ;
      RECT 879.475000 0.000000 881.325000 0.630000 ;
      RECT 877.200000 0.000000 879.055000 0.630000 ;
      RECT 874.930000 0.000000 876.780000 0.630000 ;
      RECT 872.660000 0.000000 874.510000 0.630000 ;
      RECT 870.385000 0.000000 872.240000 0.630000 ;
      RECT 868.115000 0.000000 869.965000 0.630000 ;
      RECT 865.840000 0.000000 867.695000 0.630000 ;
      RECT 863.570000 0.000000 865.420000 0.630000 ;
      RECT 861.300000 0.000000 863.150000 0.630000 ;
      RECT 859.025000 0.000000 860.880000 0.630000 ;
      RECT 856.755000 0.000000 858.605000 0.630000 ;
      RECT 854.480000 0.000000 856.335000 0.630000 ;
      RECT 852.210000 0.000000 854.060000 0.630000 ;
      RECT 849.940000 0.000000 851.790000 0.630000 ;
      RECT 847.665000 0.000000 849.520000 0.630000 ;
      RECT 845.395000 0.000000 847.245000 0.630000 ;
      RECT 843.120000 0.000000 844.975000 0.630000 ;
      RECT 840.850000 0.000000 842.700000 0.630000 ;
      RECT 838.580000 0.000000 840.430000 0.630000 ;
      RECT 836.305000 0.000000 838.160000 0.630000 ;
      RECT 834.035000 0.000000 835.885000 0.630000 ;
      RECT 831.760000 0.000000 833.615000 0.630000 ;
      RECT 829.490000 0.000000 831.340000 0.630000 ;
      RECT 827.220000 0.000000 829.070000 0.630000 ;
      RECT 824.945000 0.000000 826.800000 0.630000 ;
      RECT 822.675000 0.000000 824.525000 0.630000 ;
      RECT 820.400000 0.000000 822.255000 0.630000 ;
      RECT 818.130000 0.000000 819.980000 0.630000 ;
      RECT 815.860000 0.000000 817.710000 0.630000 ;
      RECT 813.585000 0.000000 815.440000 0.630000 ;
      RECT 811.315000 0.000000 813.165000 0.630000 ;
      RECT 809.040000 0.000000 810.895000 0.630000 ;
      RECT 806.770000 0.000000 808.620000 0.630000 ;
      RECT 804.500000 0.000000 806.350000 0.630000 ;
      RECT 802.225000 0.000000 804.080000 0.630000 ;
      RECT 799.955000 0.000000 801.805000 0.630000 ;
      RECT 797.680000 0.000000 799.535000 0.630000 ;
      RECT 795.410000 0.000000 797.260000 0.630000 ;
      RECT 793.140000 0.000000 794.990000 0.630000 ;
      RECT 790.865000 0.000000 792.720000 0.630000 ;
      RECT 788.595000 0.000000 790.445000 0.630000 ;
      RECT 786.320000 0.000000 788.175000 0.630000 ;
      RECT 784.050000 0.000000 785.900000 0.630000 ;
      RECT 781.780000 0.000000 783.630000 0.630000 ;
      RECT 779.505000 0.000000 781.360000 0.630000 ;
      RECT 777.235000 0.000000 779.085000 0.630000 ;
      RECT 774.960000 0.000000 776.815000 0.630000 ;
      RECT 772.690000 0.000000 774.540000 0.630000 ;
      RECT 770.420000 0.000000 772.270000 0.630000 ;
      RECT 768.145000 0.000000 770.000000 0.630000 ;
      RECT 765.875000 0.000000 767.725000 0.630000 ;
      RECT 763.600000 0.000000 765.455000 0.630000 ;
      RECT 761.330000 0.000000 763.180000 0.630000 ;
      RECT 759.060000 0.000000 760.910000 0.630000 ;
      RECT 756.785000 0.000000 758.640000 0.630000 ;
      RECT 754.515000 0.000000 756.365000 0.630000 ;
      RECT 752.240000 0.000000 754.095000 0.630000 ;
      RECT 749.970000 0.000000 751.820000 0.630000 ;
      RECT 747.700000 0.000000 749.550000 0.630000 ;
      RECT 745.425000 0.000000 747.280000 0.630000 ;
      RECT 743.155000 0.000000 745.005000 0.630000 ;
      RECT 740.880000 0.000000 742.735000 0.630000 ;
      RECT 738.610000 0.000000 740.460000 0.630000 ;
      RECT 736.340000 0.000000 738.190000 0.630000 ;
      RECT 734.065000 0.000000 735.920000 0.630000 ;
      RECT 731.795000 0.000000 733.645000 0.630000 ;
      RECT 729.520000 0.000000 731.375000 0.630000 ;
      RECT 727.250000 0.000000 729.100000 0.630000 ;
      RECT 724.980000 0.000000 726.830000 0.630000 ;
      RECT 722.705000 0.000000 724.560000 0.630000 ;
      RECT 720.435000 0.000000 722.285000 0.630000 ;
      RECT 718.160000 0.000000 720.015000 0.630000 ;
      RECT 715.890000 0.000000 717.740000 0.630000 ;
      RECT 713.620000 0.000000 715.470000 0.630000 ;
      RECT 711.345000 0.000000 713.200000 0.630000 ;
      RECT 709.075000 0.000000 710.925000 0.630000 ;
      RECT 706.800000 0.000000 708.655000 0.630000 ;
      RECT 704.530000 0.000000 706.380000 0.630000 ;
      RECT 702.260000 0.000000 704.110000 0.630000 ;
      RECT 699.985000 0.000000 701.840000 0.630000 ;
      RECT 697.715000 0.000000 699.565000 0.630000 ;
      RECT 695.440000 0.000000 697.295000 0.630000 ;
      RECT 693.170000 0.000000 695.020000 0.630000 ;
      RECT 690.900000 0.000000 692.750000 0.630000 ;
      RECT 688.625000 0.000000 690.480000 0.630000 ;
      RECT 686.355000 0.000000 688.205000 0.630000 ;
      RECT 684.080000 0.000000 685.935000 0.630000 ;
      RECT 681.810000 0.000000 683.660000 0.630000 ;
      RECT 679.540000 0.000000 681.390000 0.630000 ;
      RECT 677.265000 0.000000 679.120000 0.630000 ;
      RECT 674.995000 0.000000 676.845000 0.630000 ;
      RECT 672.720000 0.000000 674.575000 0.630000 ;
      RECT 670.450000 0.000000 672.300000 0.630000 ;
      RECT 668.180000 0.000000 670.030000 0.630000 ;
      RECT 665.905000 0.000000 667.760000 0.630000 ;
      RECT 663.635000 0.000000 665.485000 0.630000 ;
      RECT 661.360000 0.000000 663.215000 0.630000 ;
      RECT 659.090000 0.000000 660.940000 0.630000 ;
      RECT 656.820000 0.000000 658.670000 0.630000 ;
      RECT 654.545000 0.000000 656.400000 0.630000 ;
      RECT 652.275000 0.000000 654.125000 0.630000 ;
      RECT 650.000000 0.000000 651.855000 0.630000 ;
      RECT 647.730000 0.000000 649.580000 0.630000 ;
      RECT 645.460000 0.000000 647.310000 0.630000 ;
      RECT 643.185000 0.000000 645.040000 0.630000 ;
      RECT 640.915000 0.000000 642.765000 0.630000 ;
      RECT 638.640000 0.000000 640.495000 0.630000 ;
      RECT 636.370000 0.000000 638.220000 0.630000 ;
      RECT 634.100000 0.000000 635.950000 0.630000 ;
      RECT 631.825000 0.000000 633.680000 0.630000 ;
      RECT 629.555000 0.000000 631.405000 0.630000 ;
      RECT 627.280000 0.000000 629.135000 0.630000 ;
      RECT 625.010000 0.000000 626.860000 0.630000 ;
      RECT 622.740000 0.000000 624.590000 0.630000 ;
      RECT 620.465000 0.000000 622.320000 0.630000 ;
      RECT 618.195000 0.000000 620.045000 0.630000 ;
      RECT 615.920000 0.000000 617.775000 0.630000 ;
      RECT 613.650000 0.000000 615.500000 0.630000 ;
      RECT 611.380000 0.000000 613.230000 0.630000 ;
      RECT 609.105000 0.000000 610.960000 0.630000 ;
      RECT 606.835000 0.000000 608.685000 0.630000 ;
      RECT 604.560000 0.000000 606.415000 0.630000 ;
      RECT 602.290000 0.000000 604.140000 0.630000 ;
      RECT 600.020000 0.000000 601.870000 0.630000 ;
      RECT 597.745000 0.000000 599.600000 0.630000 ;
      RECT 595.475000 0.000000 597.325000 0.630000 ;
      RECT 593.200000 0.000000 595.055000 0.630000 ;
      RECT 590.930000 0.000000 592.780000 0.630000 ;
      RECT 588.660000 0.000000 590.510000 0.630000 ;
      RECT 586.385000 0.000000 588.240000 0.630000 ;
      RECT 584.115000 0.000000 585.965000 0.630000 ;
      RECT 581.840000 0.000000 583.695000 0.630000 ;
      RECT 579.570000 0.000000 581.420000 0.630000 ;
      RECT 577.300000 0.000000 579.150000 0.630000 ;
      RECT 575.025000 0.000000 576.880000 0.630000 ;
      RECT 572.755000 0.000000 574.605000 0.630000 ;
      RECT 570.480000 0.000000 572.335000 0.630000 ;
      RECT 568.210000 0.000000 570.060000 0.630000 ;
      RECT 565.940000 0.000000 567.790000 0.630000 ;
      RECT 563.665000 0.000000 565.520000 0.630000 ;
      RECT 561.395000 0.000000 563.245000 0.630000 ;
      RECT 559.120000 0.000000 560.975000 0.630000 ;
      RECT 556.850000 0.000000 558.700000 0.630000 ;
      RECT 554.580000 0.000000 556.430000 0.630000 ;
      RECT 552.305000 0.000000 554.160000 0.630000 ;
      RECT 550.035000 0.000000 551.885000 0.630000 ;
      RECT 547.760000 0.000000 549.615000 0.630000 ;
      RECT 545.490000 0.000000 547.340000 0.630000 ;
      RECT 543.220000 0.000000 545.070000 0.630000 ;
      RECT 540.945000 0.000000 542.800000 0.630000 ;
      RECT 538.675000 0.000000 540.525000 0.630000 ;
      RECT 536.400000 0.000000 538.255000 0.630000 ;
      RECT 534.130000 0.000000 535.980000 0.630000 ;
      RECT 531.860000 0.000000 533.710000 0.630000 ;
      RECT 529.585000 0.000000 531.440000 0.630000 ;
      RECT 527.315000 0.000000 529.165000 0.630000 ;
      RECT 525.040000 0.000000 526.895000 0.630000 ;
      RECT 522.770000 0.000000 524.620000 0.630000 ;
      RECT 520.500000 0.000000 522.350000 0.630000 ;
      RECT 518.225000 0.000000 520.080000 0.630000 ;
      RECT 515.955000 0.000000 517.805000 0.630000 ;
      RECT 513.680000 0.000000 515.535000 0.630000 ;
      RECT 511.410000 0.000000 513.260000 0.630000 ;
      RECT 509.140000 0.000000 510.990000 0.630000 ;
      RECT 506.865000 0.000000 508.720000 0.630000 ;
      RECT 504.595000 0.000000 506.445000 0.630000 ;
      RECT 502.320000 0.000000 504.175000 0.630000 ;
      RECT 500.050000 0.000000 501.900000 0.630000 ;
      RECT 497.780000 0.000000 499.630000 0.630000 ;
      RECT 495.505000 0.000000 497.360000 0.630000 ;
      RECT 493.235000 0.000000 495.085000 0.630000 ;
      RECT 490.960000 0.000000 492.815000 0.630000 ;
      RECT 488.690000 0.000000 490.540000 0.630000 ;
      RECT 486.420000 0.000000 488.270000 0.630000 ;
      RECT 484.145000 0.000000 486.000000 0.630000 ;
      RECT 481.875000 0.000000 483.725000 0.630000 ;
      RECT 479.600000 0.000000 481.455000 0.630000 ;
      RECT 477.330000 0.000000 479.180000 0.630000 ;
      RECT 475.060000 0.000000 476.910000 0.630000 ;
      RECT 472.785000 0.000000 474.640000 0.630000 ;
      RECT 470.515000 0.000000 472.365000 0.630000 ;
      RECT 468.240000 0.000000 470.095000 0.630000 ;
      RECT 465.970000 0.000000 467.820000 0.630000 ;
      RECT 463.700000 0.000000 465.550000 0.630000 ;
      RECT 461.425000 0.000000 463.280000 0.630000 ;
      RECT 459.155000 0.000000 461.005000 0.630000 ;
      RECT 456.880000 0.000000 458.735000 0.630000 ;
      RECT 454.610000 0.000000 456.460000 0.630000 ;
      RECT 452.340000 0.000000 454.190000 0.630000 ;
      RECT 450.065000 0.000000 451.920000 0.630000 ;
      RECT 447.795000 0.000000 449.645000 0.630000 ;
      RECT 445.520000 0.000000 447.375000 0.630000 ;
      RECT 443.250000 0.000000 445.100000 0.630000 ;
      RECT 440.980000 0.000000 442.830000 0.630000 ;
      RECT 438.705000 0.000000 440.560000 0.630000 ;
      RECT 436.435000 0.000000 438.285000 0.630000 ;
      RECT 434.160000 0.000000 436.015000 0.630000 ;
      RECT 431.890000 0.000000 433.740000 0.630000 ;
      RECT 429.620000 0.000000 431.470000 0.630000 ;
      RECT 427.345000 0.000000 429.200000 0.630000 ;
      RECT 425.075000 0.000000 426.925000 0.630000 ;
      RECT 422.800000 0.000000 424.655000 0.630000 ;
      RECT 420.530000 0.000000 422.380000 0.630000 ;
      RECT 418.260000 0.000000 420.110000 0.630000 ;
      RECT 415.985000 0.000000 417.840000 0.630000 ;
      RECT 413.715000 0.000000 415.565000 0.630000 ;
      RECT 411.440000 0.000000 413.295000 0.630000 ;
      RECT 409.170000 0.000000 411.020000 0.630000 ;
      RECT 406.900000 0.000000 408.750000 0.630000 ;
      RECT 404.625000 0.000000 406.480000 0.630000 ;
      RECT 402.355000 0.000000 404.205000 0.630000 ;
      RECT 400.080000 0.000000 401.935000 0.630000 ;
      RECT 397.810000 0.000000 399.660000 0.630000 ;
      RECT 395.540000 0.000000 397.390000 0.630000 ;
      RECT 393.265000 0.000000 395.120000 0.630000 ;
      RECT 390.995000 0.000000 392.845000 0.630000 ;
      RECT 388.720000 0.000000 390.575000 0.630000 ;
      RECT 386.450000 0.000000 388.300000 0.630000 ;
      RECT 384.180000 0.000000 386.030000 0.630000 ;
      RECT 381.905000 0.000000 383.760000 0.630000 ;
      RECT 379.635000 0.000000 381.485000 0.630000 ;
      RECT 377.360000 0.000000 379.215000 0.630000 ;
      RECT 375.090000 0.000000 376.940000 0.630000 ;
      RECT 372.820000 0.000000 374.670000 0.630000 ;
      RECT 370.545000 0.000000 372.400000 0.630000 ;
      RECT 368.275000 0.000000 370.125000 0.630000 ;
      RECT 366.000000 0.000000 367.855000 0.630000 ;
      RECT 363.730000 0.000000 365.580000 0.630000 ;
      RECT 361.460000 0.000000 363.310000 0.630000 ;
      RECT 359.185000 0.000000 361.040000 0.630000 ;
      RECT 356.915000 0.000000 358.765000 0.630000 ;
      RECT 354.640000 0.000000 356.495000 0.630000 ;
      RECT 352.370000 0.000000 354.220000 0.630000 ;
      RECT 350.100000 0.000000 351.950000 0.630000 ;
      RECT 347.825000 0.000000 349.680000 0.630000 ;
      RECT 345.555000 0.000000 347.405000 0.630000 ;
      RECT 343.280000 0.000000 345.135000 0.630000 ;
      RECT 341.010000 0.000000 342.860000 0.630000 ;
      RECT 338.740000 0.000000 340.590000 0.630000 ;
      RECT 336.465000 0.000000 338.320000 0.630000 ;
      RECT 334.195000 0.000000 336.045000 0.630000 ;
      RECT 331.920000 0.000000 333.775000 0.630000 ;
      RECT 329.650000 0.000000 331.500000 0.630000 ;
      RECT 327.380000 0.000000 329.230000 0.630000 ;
      RECT 325.105000 0.000000 326.960000 0.630000 ;
      RECT 322.835000 0.000000 324.685000 0.630000 ;
      RECT 320.560000 0.000000 322.415000 0.630000 ;
      RECT 318.290000 0.000000 320.140000 0.630000 ;
      RECT 316.020000 0.000000 317.870000 0.630000 ;
      RECT 313.745000 0.000000 315.600000 0.630000 ;
      RECT 311.475000 0.000000 313.325000 0.630000 ;
      RECT 309.200000 0.000000 311.055000 0.630000 ;
      RECT 306.930000 0.000000 308.780000 0.630000 ;
      RECT 304.660000 0.000000 306.510000 0.630000 ;
      RECT 302.385000 0.000000 304.240000 0.630000 ;
      RECT 300.115000 0.000000 301.965000 0.630000 ;
      RECT 297.840000 0.000000 299.695000 0.630000 ;
      RECT 295.570000 0.000000 297.420000 0.630000 ;
      RECT 293.300000 0.000000 295.150000 0.630000 ;
      RECT 291.025000 0.000000 292.880000 0.630000 ;
      RECT 288.755000 0.000000 290.605000 0.630000 ;
      RECT 286.480000 0.000000 288.335000 0.630000 ;
      RECT 284.210000 0.000000 286.060000 0.630000 ;
      RECT 281.940000 0.000000 283.790000 0.630000 ;
      RECT 279.665000 0.000000 281.520000 0.630000 ;
      RECT 277.395000 0.000000 279.245000 0.630000 ;
      RECT 275.120000 0.000000 276.975000 0.630000 ;
      RECT 272.850000 0.000000 274.700000 0.630000 ;
      RECT 270.580000 0.000000 272.430000 0.630000 ;
      RECT 268.305000 0.000000 270.160000 0.630000 ;
      RECT 266.035000 0.000000 267.885000 0.630000 ;
      RECT 263.760000 0.000000 265.615000 0.630000 ;
      RECT 261.490000 0.000000 263.340000 0.630000 ;
      RECT 259.220000 0.000000 261.070000 0.630000 ;
      RECT 256.945000 0.000000 258.800000 0.630000 ;
      RECT 254.675000 0.000000 256.525000 0.630000 ;
      RECT 252.400000 0.000000 254.255000 0.630000 ;
      RECT 250.130000 0.000000 251.980000 0.630000 ;
      RECT 247.860000 0.000000 249.710000 0.630000 ;
      RECT 245.585000 0.000000 247.440000 0.630000 ;
      RECT 243.315000 0.000000 245.165000 0.630000 ;
      RECT 241.040000 0.000000 242.895000 0.630000 ;
      RECT 238.770000 0.000000 240.620000 0.630000 ;
      RECT 236.500000 0.000000 238.350000 0.630000 ;
      RECT 234.225000 0.000000 236.080000 0.630000 ;
      RECT 231.955000 0.000000 233.805000 0.630000 ;
      RECT 229.680000 0.000000 231.535000 0.630000 ;
      RECT 227.410000 0.000000 229.260000 0.630000 ;
      RECT 225.140000 0.000000 226.990000 0.630000 ;
      RECT 222.865000 0.000000 224.720000 0.630000 ;
      RECT 220.595000 0.000000 222.445000 0.630000 ;
      RECT 218.320000 0.000000 220.175000 0.630000 ;
      RECT 216.050000 0.000000 217.900000 0.630000 ;
      RECT 213.780000 0.000000 215.630000 0.630000 ;
      RECT 211.505000 0.000000 213.360000 0.630000 ;
      RECT 209.235000 0.000000 211.085000 0.630000 ;
      RECT 206.960000 0.000000 208.815000 0.630000 ;
      RECT 204.690000 0.000000 206.540000 0.630000 ;
      RECT 202.420000 0.000000 204.270000 0.630000 ;
      RECT 200.145000 0.000000 202.000000 0.630000 ;
      RECT 197.875000 0.000000 199.725000 0.630000 ;
      RECT 195.600000 0.000000 197.455000 0.630000 ;
      RECT 193.330000 0.000000 195.180000 0.630000 ;
      RECT 191.060000 0.000000 192.910000 0.630000 ;
      RECT 188.785000 0.000000 190.640000 0.630000 ;
      RECT 186.515000 0.000000 188.365000 0.630000 ;
      RECT 184.240000 0.000000 186.095000 0.630000 ;
      RECT 181.970000 0.000000 183.820000 0.630000 ;
      RECT 179.700000 0.000000 181.550000 0.630000 ;
      RECT 177.425000 0.000000 179.280000 0.630000 ;
      RECT 175.155000 0.000000 177.005000 0.630000 ;
      RECT 172.880000 0.000000 174.735000 0.630000 ;
      RECT 170.610000 0.000000 172.460000 0.630000 ;
      RECT 168.340000 0.000000 170.190000 0.630000 ;
      RECT 166.065000 0.000000 167.920000 0.630000 ;
      RECT 163.795000 0.000000 165.645000 0.630000 ;
      RECT 161.520000 0.000000 163.375000 0.630000 ;
      RECT 159.250000 0.000000 161.100000 0.630000 ;
      RECT 156.980000 0.000000 158.830000 0.630000 ;
      RECT 154.705000 0.000000 156.560000 0.630000 ;
      RECT 152.435000 0.000000 154.285000 0.630000 ;
      RECT 150.160000 0.000000 152.015000 0.630000 ;
      RECT 147.890000 0.000000 149.740000 0.630000 ;
      RECT 145.620000 0.000000 147.470000 0.630000 ;
      RECT 143.345000 0.000000 145.200000 0.630000 ;
      RECT 141.075000 0.000000 142.925000 0.630000 ;
      RECT 138.800000 0.000000 140.655000 0.630000 ;
      RECT 136.530000 0.000000 138.380000 0.630000 ;
      RECT 134.260000 0.000000 136.110000 0.630000 ;
      RECT 131.985000 0.000000 133.840000 0.630000 ;
      RECT 129.715000 0.000000 131.565000 0.630000 ;
      RECT 127.440000 0.000000 129.295000 0.630000 ;
      RECT 125.170000 0.000000 127.020000 0.630000 ;
      RECT 122.900000 0.000000 124.750000 0.630000 ;
      RECT 120.625000 0.000000 122.480000 0.630000 ;
      RECT 118.355000 0.000000 120.205000 0.630000 ;
      RECT 116.080000 0.000000 117.935000 0.630000 ;
      RECT 113.810000 0.000000 115.660000 0.630000 ;
      RECT 111.540000 0.000000 113.390000 0.630000 ;
      RECT 109.265000 0.000000 111.120000 0.630000 ;
      RECT 106.995000 0.000000 108.845000 0.630000 ;
      RECT 104.720000 0.000000 106.575000 0.630000 ;
      RECT 102.450000 0.000000 104.300000 0.630000 ;
      RECT 100.180000 0.000000 102.030000 0.630000 ;
      RECT 97.905000 0.000000 99.760000 0.630000 ;
      RECT 95.635000 0.000000 97.485000 0.630000 ;
      RECT 93.360000 0.000000 95.215000 0.630000 ;
      RECT 91.090000 0.000000 92.940000 0.630000 ;
      RECT 88.820000 0.000000 90.670000 0.630000 ;
      RECT 86.545000 0.000000 88.400000 0.630000 ;
      RECT 84.275000 0.000000 86.125000 0.630000 ;
      RECT 82.000000 0.000000 83.855000 0.630000 ;
      RECT 79.730000 0.000000 81.580000 0.630000 ;
      RECT 77.460000 0.000000 79.310000 0.630000 ;
      RECT 75.185000 0.000000 77.040000 0.630000 ;
      RECT 72.915000 0.000000 74.765000 0.630000 ;
      RECT 70.640000 0.000000 72.495000 0.630000 ;
      RECT 68.370000 0.000000 70.220000 0.630000 ;
      RECT 66.100000 0.000000 67.950000 0.630000 ;
      RECT 63.825000 0.000000 65.680000 0.630000 ;
      RECT 61.555000 0.000000 63.405000 0.630000 ;
      RECT 59.280000 0.000000 61.135000 0.630000 ;
      RECT 57.010000 0.000000 58.860000 0.630000 ;
      RECT 54.740000 0.000000 56.590000 0.630000 ;
      RECT 52.465000 0.000000 54.320000 0.630000 ;
      RECT 50.195000 0.000000 52.045000 0.630000 ;
      RECT 47.920000 0.000000 49.775000 0.630000 ;
      RECT 45.650000 0.000000 47.500000 0.630000 ;
      RECT 43.380000 0.000000 45.230000 0.630000 ;
      RECT 41.105000 0.000000 42.960000 0.630000 ;
      RECT 38.835000 0.000000 40.685000 0.630000 ;
      RECT 36.560000 0.000000 38.415000 0.630000 ;
      RECT 34.290000 0.000000 36.140000 0.630000 ;
      RECT 32.020000 0.000000 33.870000 0.630000 ;
      RECT 29.745000 0.000000 31.600000 0.630000 ;
      RECT 27.475000 0.000000 29.325000 0.630000 ;
      RECT 25.200000 0.000000 27.055000 0.630000 ;
      RECT 22.930000 0.000000 24.780000 0.630000 ;
      RECT 20.660000 0.000000 22.510000 0.630000 ;
      RECT 18.385000 0.000000 20.240000 0.630000 ;
      RECT 16.115000 0.000000 17.965000 0.630000 ;
      RECT 13.840000 0.000000 15.695000 0.630000 ;
      RECT 11.570000 0.000000 13.420000 0.630000 ;
      RECT 9.300000 0.000000 11.150000 0.630000 ;
      RECT 7.025000 0.000000 8.880000 0.630000 ;
      RECT 4.755000 0.000000 6.605000 0.630000 ;
      RECT 2.480000 0.000000 4.335000 0.630000 ;
      RECT 1.820000 0.000000 2.060000 0.630000 ;
      RECT 0.000000 0.000000 1.400000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 916.940000 1120.100000 919.700000 ;
      RECT 1.100000 916.330000 1120.100000 916.940000 ;
      RECT 1.100000 916.040000 1119.000000 916.330000 ;
      RECT 0.000000 915.430000 1119.000000 916.040000 ;
      RECT 0.000000 902.755000 1120.100000 915.430000 ;
      RECT 1.100000 902.435000 1120.100000 902.755000 ;
      RECT 1.100000 901.855000 1119.000000 902.435000 ;
      RECT 0.000000 901.535000 1119.000000 901.855000 ;
      RECT 0.000000 885.400000 1120.100000 901.535000 ;
      RECT 1.100000 884.750000 1120.100000 885.400000 ;
      RECT 1.100000 884.500000 1119.000000 884.750000 ;
      RECT 0.000000 883.850000 1119.000000 884.500000 ;
      RECT 0.000000 868.050000 1120.100000 883.850000 ;
      RECT 1.100000 867.150000 1120.100000 868.050000 ;
      RECT 0.000000 867.065000 1120.100000 867.150000 ;
      RECT 0.000000 866.165000 1119.000000 867.065000 ;
      RECT 0.000000 850.700000 1120.100000 866.165000 ;
      RECT 1.100000 849.800000 1120.100000 850.700000 ;
      RECT 0.000000 849.380000 1120.100000 849.800000 ;
      RECT 0.000000 848.480000 1119.000000 849.380000 ;
      RECT 0.000000 833.345000 1120.100000 848.480000 ;
      RECT 1.100000 832.445000 1120.100000 833.345000 ;
      RECT 0.000000 831.690000 1120.100000 832.445000 ;
      RECT 0.000000 830.790000 1119.000000 831.690000 ;
      RECT 0.000000 815.995000 1120.100000 830.790000 ;
      RECT 1.100000 815.095000 1120.100000 815.995000 ;
      RECT 0.000000 814.005000 1120.100000 815.095000 ;
      RECT 0.000000 813.105000 1119.000000 814.005000 ;
      RECT 0.000000 798.640000 1120.100000 813.105000 ;
      RECT 1.100000 797.740000 1120.100000 798.640000 ;
      RECT 0.000000 796.320000 1120.100000 797.740000 ;
      RECT 0.000000 795.420000 1119.000000 796.320000 ;
      RECT 0.000000 781.290000 1120.100000 795.420000 ;
      RECT 1.100000 780.390000 1120.100000 781.290000 ;
      RECT 0.000000 778.635000 1120.100000 780.390000 ;
      RECT 0.000000 777.735000 1119.000000 778.635000 ;
      RECT 0.000000 763.940000 1120.100000 777.735000 ;
      RECT 1.100000 763.040000 1120.100000 763.940000 ;
      RECT 0.000000 760.950000 1120.100000 763.040000 ;
      RECT 0.000000 760.050000 1119.000000 760.950000 ;
      RECT 0.000000 746.585000 1120.100000 760.050000 ;
      RECT 1.100000 745.685000 1120.100000 746.585000 ;
      RECT 0.000000 743.260000 1120.100000 745.685000 ;
      RECT 0.000000 742.360000 1119.000000 743.260000 ;
      RECT 0.000000 729.235000 1120.100000 742.360000 ;
      RECT 1.100000 728.335000 1120.100000 729.235000 ;
      RECT 0.000000 725.575000 1120.100000 728.335000 ;
      RECT 0.000000 724.675000 1119.000000 725.575000 ;
      RECT 0.000000 711.880000 1120.100000 724.675000 ;
      RECT 1.100000 710.980000 1120.100000 711.880000 ;
      RECT 0.000000 707.890000 1120.100000 710.980000 ;
      RECT 0.000000 706.990000 1119.000000 707.890000 ;
      RECT 0.000000 694.530000 1120.100000 706.990000 ;
      RECT 1.100000 693.630000 1120.100000 694.530000 ;
      RECT 0.000000 690.205000 1120.100000 693.630000 ;
      RECT 0.000000 689.305000 1119.000000 690.205000 ;
      RECT 0.000000 677.180000 1120.100000 689.305000 ;
      RECT 1.100000 676.280000 1120.100000 677.180000 ;
      RECT 0.000000 672.520000 1120.100000 676.280000 ;
      RECT 0.000000 671.620000 1119.000000 672.520000 ;
      RECT 0.000000 659.825000 1120.100000 671.620000 ;
      RECT 1.100000 658.925000 1120.100000 659.825000 ;
      RECT 0.000000 654.830000 1120.100000 658.925000 ;
      RECT 0.000000 653.930000 1119.000000 654.830000 ;
      RECT 0.000000 642.475000 1120.100000 653.930000 ;
      RECT 1.100000 641.575000 1120.100000 642.475000 ;
      RECT 0.000000 637.145000 1120.100000 641.575000 ;
      RECT 0.000000 636.245000 1119.000000 637.145000 ;
      RECT 0.000000 625.120000 1120.100000 636.245000 ;
      RECT 1.100000 624.220000 1120.100000 625.120000 ;
      RECT 0.000000 619.460000 1120.100000 624.220000 ;
      RECT 0.000000 618.560000 1119.000000 619.460000 ;
      RECT 0.000000 607.770000 1120.100000 618.560000 ;
      RECT 1.100000 606.870000 1120.100000 607.770000 ;
      RECT 0.000000 601.775000 1120.100000 606.870000 ;
      RECT 0.000000 600.875000 1119.000000 601.775000 ;
      RECT 0.000000 590.420000 1120.100000 600.875000 ;
      RECT 1.100000 589.520000 1120.100000 590.420000 ;
      RECT 0.000000 584.090000 1120.100000 589.520000 ;
      RECT 0.000000 583.190000 1119.000000 584.090000 ;
      RECT 0.000000 573.065000 1120.100000 583.190000 ;
      RECT 1.100000 572.165000 1120.100000 573.065000 ;
      RECT 0.000000 566.400000 1120.100000 572.165000 ;
      RECT 0.000000 565.500000 1119.000000 566.400000 ;
      RECT 0.000000 555.715000 1120.100000 565.500000 ;
      RECT 1.100000 554.815000 1120.100000 555.715000 ;
      RECT 0.000000 548.715000 1120.100000 554.815000 ;
      RECT 0.000000 547.815000 1119.000000 548.715000 ;
      RECT 0.000000 538.360000 1120.100000 547.815000 ;
      RECT 1.100000 537.460000 1120.100000 538.360000 ;
      RECT 0.000000 531.030000 1120.100000 537.460000 ;
      RECT 0.000000 530.130000 1119.000000 531.030000 ;
      RECT 0.000000 521.010000 1120.100000 530.130000 ;
      RECT 1.100000 520.110000 1120.100000 521.010000 ;
      RECT 0.000000 513.345000 1120.100000 520.110000 ;
      RECT 0.000000 512.445000 1119.000000 513.345000 ;
      RECT 0.000000 503.660000 1120.100000 512.445000 ;
      RECT 1.100000 502.760000 1120.100000 503.660000 ;
      RECT 0.000000 495.660000 1120.100000 502.760000 ;
      RECT 0.000000 494.760000 1119.000000 495.660000 ;
      RECT 0.000000 486.305000 1120.100000 494.760000 ;
      RECT 1.100000 485.405000 1120.100000 486.305000 ;
      RECT 0.000000 477.970000 1120.100000 485.405000 ;
      RECT 0.000000 477.070000 1119.000000 477.970000 ;
      RECT 0.000000 468.955000 1120.100000 477.070000 ;
      RECT 1.100000 468.055000 1120.100000 468.955000 ;
      RECT 0.000000 460.285000 1120.100000 468.055000 ;
      RECT 0.000000 459.385000 1119.000000 460.285000 ;
      RECT 0.000000 451.600000 1120.100000 459.385000 ;
      RECT 1.100000 450.700000 1120.100000 451.600000 ;
      RECT 0.000000 442.600000 1120.100000 450.700000 ;
      RECT 0.000000 441.700000 1119.000000 442.600000 ;
      RECT 0.000000 434.250000 1120.100000 441.700000 ;
      RECT 1.100000 433.350000 1120.100000 434.250000 ;
      RECT 0.000000 424.915000 1120.100000 433.350000 ;
      RECT 0.000000 424.015000 1119.000000 424.915000 ;
      RECT 0.000000 416.900000 1120.100000 424.015000 ;
      RECT 1.100000 416.000000 1120.100000 416.900000 ;
      RECT 0.000000 407.230000 1120.100000 416.000000 ;
      RECT 0.000000 406.330000 1119.000000 407.230000 ;
      RECT 0.000000 399.545000 1120.100000 406.330000 ;
      RECT 1.100000 398.645000 1120.100000 399.545000 ;
      RECT 0.000000 389.540000 1120.100000 398.645000 ;
      RECT 0.000000 388.640000 1119.000000 389.540000 ;
      RECT 0.000000 382.195000 1120.100000 388.640000 ;
      RECT 1.100000 381.295000 1120.100000 382.195000 ;
      RECT 0.000000 371.855000 1120.100000 381.295000 ;
      RECT 0.000000 370.955000 1119.000000 371.855000 ;
      RECT 0.000000 364.840000 1120.100000 370.955000 ;
      RECT 1.100000 363.940000 1120.100000 364.840000 ;
      RECT 0.000000 354.170000 1120.100000 363.940000 ;
      RECT 0.000000 353.270000 1119.000000 354.170000 ;
      RECT 0.000000 347.490000 1120.100000 353.270000 ;
      RECT 1.100000 346.590000 1120.100000 347.490000 ;
      RECT 0.000000 336.485000 1120.100000 346.590000 ;
      RECT 0.000000 335.585000 1119.000000 336.485000 ;
      RECT 0.000000 330.140000 1120.100000 335.585000 ;
      RECT 1.100000 329.240000 1120.100000 330.140000 ;
      RECT 0.000000 318.800000 1120.100000 329.240000 ;
      RECT 0.000000 317.900000 1119.000000 318.800000 ;
      RECT 0.000000 312.785000 1120.100000 317.900000 ;
      RECT 1.100000 311.885000 1120.100000 312.785000 ;
      RECT 0.000000 301.110000 1120.100000 311.885000 ;
      RECT 0.000000 300.210000 1119.000000 301.110000 ;
      RECT 0.000000 295.435000 1120.100000 300.210000 ;
      RECT 1.100000 294.535000 1120.100000 295.435000 ;
      RECT 0.000000 283.425000 1120.100000 294.535000 ;
      RECT 0.000000 282.525000 1119.000000 283.425000 ;
      RECT 0.000000 278.080000 1120.100000 282.525000 ;
      RECT 1.100000 277.180000 1120.100000 278.080000 ;
      RECT 0.000000 265.740000 1120.100000 277.180000 ;
      RECT 0.000000 264.840000 1119.000000 265.740000 ;
      RECT 0.000000 260.730000 1120.100000 264.840000 ;
      RECT 1.100000 259.830000 1120.100000 260.730000 ;
      RECT 0.000000 248.055000 1120.100000 259.830000 ;
      RECT 0.000000 247.155000 1119.000000 248.055000 ;
      RECT 0.000000 243.380000 1120.100000 247.155000 ;
      RECT 1.100000 242.480000 1120.100000 243.380000 ;
      RECT 0.000000 230.370000 1120.100000 242.480000 ;
      RECT 0.000000 229.470000 1119.000000 230.370000 ;
      RECT 0.000000 226.025000 1120.100000 229.470000 ;
      RECT 1.100000 225.125000 1120.100000 226.025000 ;
      RECT 0.000000 212.680000 1120.100000 225.125000 ;
      RECT 0.000000 211.780000 1119.000000 212.680000 ;
      RECT 0.000000 208.675000 1120.100000 211.780000 ;
      RECT 1.100000 207.775000 1120.100000 208.675000 ;
      RECT 0.000000 194.995000 1120.100000 207.775000 ;
      RECT 0.000000 194.095000 1119.000000 194.995000 ;
      RECT 0.000000 191.320000 1120.100000 194.095000 ;
      RECT 1.100000 190.420000 1120.100000 191.320000 ;
      RECT 0.000000 177.310000 1120.100000 190.420000 ;
      RECT 0.000000 176.410000 1119.000000 177.310000 ;
      RECT 0.000000 173.970000 1120.100000 176.410000 ;
      RECT 1.100000 173.070000 1120.100000 173.970000 ;
      RECT 0.000000 159.625000 1120.100000 173.070000 ;
      RECT 0.000000 158.725000 1119.000000 159.625000 ;
      RECT 0.000000 156.620000 1120.100000 158.725000 ;
      RECT 1.100000 155.720000 1120.100000 156.620000 ;
      RECT 0.000000 141.940000 1120.100000 155.720000 ;
      RECT 0.000000 141.040000 1119.000000 141.940000 ;
      RECT 0.000000 139.265000 1120.100000 141.040000 ;
      RECT 1.100000 138.365000 1120.100000 139.265000 ;
      RECT 0.000000 124.250000 1120.100000 138.365000 ;
      RECT 0.000000 123.350000 1119.000000 124.250000 ;
      RECT 0.000000 121.915000 1120.100000 123.350000 ;
      RECT 1.100000 121.015000 1120.100000 121.915000 ;
      RECT 0.000000 106.565000 1120.100000 121.015000 ;
      RECT 0.000000 105.665000 1119.000000 106.565000 ;
      RECT 0.000000 104.560000 1120.100000 105.665000 ;
      RECT 1.100000 103.660000 1120.100000 104.560000 ;
      RECT 0.000000 88.880000 1120.100000 103.660000 ;
      RECT 0.000000 87.980000 1119.000000 88.880000 ;
      RECT 0.000000 87.210000 1120.100000 87.980000 ;
      RECT 1.100000 86.310000 1120.100000 87.210000 ;
      RECT 0.000000 71.195000 1120.100000 86.310000 ;
      RECT 0.000000 70.295000 1119.000000 71.195000 ;
      RECT 0.000000 69.860000 1120.100000 70.295000 ;
      RECT 1.100000 68.960000 1120.100000 69.860000 ;
      RECT 0.000000 53.510000 1120.100000 68.960000 ;
      RECT 0.000000 52.610000 1119.000000 53.510000 ;
      RECT 0.000000 52.505000 1120.100000 52.610000 ;
      RECT 1.100000 51.605000 1120.100000 52.505000 ;
      RECT 0.000000 35.820000 1120.100000 51.605000 ;
      RECT 0.000000 35.155000 1119.000000 35.820000 ;
      RECT 1.100000 34.920000 1119.000000 35.155000 ;
      RECT 1.100000 34.255000 1120.100000 34.920000 ;
      RECT 0.000000 18.135000 1120.100000 34.255000 ;
      RECT 0.000000 17.800000 1119.000000 18.135000 ;
      RECT 1.100000 17.235000 1119.000000 17.800000 ;
      RECT 1.100000 16.900000 1120.100000 17.235000 ;
      RECT 0.000000 3.770000 1120.100000 16.900000 ;
      RECT 1.100000 3.160000 1120.100000 3.770000 ;
      RECT 1.100000 2.870000 1119.000000 3.160000 ;
      RECT 0.000000 2.260000 1119.000000 2.870000 ;
      RECT 0.000000 0.000000 1120.100000 2.260000 ;
    LAYER met4 ;
      RECT 0.000000 916.880000 1120.100000 919.700000 ;
      RECT 4.360000 912.880000 1115.740000 916.880000 ;
      RECT 1114.340000 5.630000 1115.740000 912.880000 ;
      RECT 8.360000 5.630000 1111.740000 912.880000 ;
      RECT 4.360000 5.630000 5.760000 912.880000 ;
      RECT 1118.340000 1.630000 1120.100000 916.880000 ;
      RECT 4.360000 1.630000 1115.740000 5.630000 ;
      RECT 0.000000 1.630000 1.760000 916.880000 ;
      RECT 0.000000 0.000000 1120.100000 1.630000 ;
  END
END user_proj_example

END LIBRARY
