##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Thu Jun 17 19:47:38 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 2820.260000 BY 3219.800000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.540000 0.000000 1.680000 0.600000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.650000 0.000000 5.790000 0.600000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.810000 0.000000 594.950000 0.600000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.130000 0.000000 200.270000 0.600000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.530000 0.000000 600.670000 0.600000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 589.090000 0.000000 589.230000 0.600000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 583.370000 0.000000 583.510000 0.600000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 577.650000 0.000000 577.790000 0.600000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.930000 0.000000 572.070000 0.600000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 383.170000 0.000000 383.310000 0.600000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 377.450000 0.000000 377.590000 0.600000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 371.730000 0.000000 371.870000 0.600000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.010000 0.000000 366.150000 0.600000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.290000 0.000000 360.430000 0.600000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 354.570000 0.000000 354.710000 0.600000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 348.850000 0.000000 348.990000 0.600000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 343.130000 0.000000 343.270000 0.600000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 337.410000 0.000000 337.550000 0.600000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.690000 0.000000 331.830000 0.600000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 325.970000 0.000000 326.110000 0.600000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 320.250000 0.000000 320.390000 0.600000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 314.530000 0.000000 314.670000 0.600000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 308.810000 0.000000 308.950000 0.600000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.090000 0.000000 303.230000 0.600000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 297.370000 0.000000 297.510000 0.600000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 291.650000 0.000000 291.790000 0.600000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 285.930000 0.000000 286.070000 0.600000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.210000 0.000000 280.350000 0.600000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.490000 0.000000 274.630000 0.600000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.770000 0.000000 268.910000 0.600000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 263.050000 0.000000 263.190000 0.600000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 257.330000 0.000000 257.470000 0.600000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 251.610000 0.000000 251.750000 0.600000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 245.890000 0.000000 246.030000 0.600000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.170000 0.000000 240.310000 0.600000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.450000 0.000000 234.590000 0.600000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.730000 0.000000 228.870000 0.600000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 223.010000 0.000000 223.150000 0.600000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 217.290000 0.000000 217.430000 0.600000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 211.570000 0.000000 211.710000 0.600000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 205.850000 0.000000 205.990000 0.600000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 194.410000 0.000000 194.550000 0.600000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 188.690000 0.000000 188.830000 0.600000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 182.970000 0.000000 183.110000 0.600000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 177.250000 0.000000 177.390000 0.600000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 171.530000 0.000000 171.670000 0.600000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 165.810000 0.000000 165.950000 0.600000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 160.090000 0.000000 160.230000 0.600000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 154.370000 0.000000 154.510000 0.600000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 148.650000 0.000000 148.790000 0.600000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 142.930000 0.000000 143.070000 0.600000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 137.210000 0.000000 137.350000 0.600000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 131.490000 0.000000 131.630000 0.600000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 125.770000 0.000000 125.910000 0.600000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 120.050000 0.000000 120.190000 0.600000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 114.330000 0.000000 114.470000 0.600000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 108.610000 0.000000 108.750000 0.600000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 102.890000 0.000000 103.030000 0.600000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 97.170000 0.000000 97.310000 0.600000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 91.450000 0.000000 91.590000 0.600000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 85.730000 0.000000 85.870000 0.600000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 80.010000 0.000000 80.150000 0.600000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.290000 0.000000 74.430000 0.600000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 68.570000 0.000000 68.710000 0.600000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.850000 0.000000 62.990000 0.600000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 57.130000 0.000000 57.270000 0.600000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 51.410000 0.000000 51.550000 0.600000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 45.690000 0.000000 45.830000 0.600000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 39.970000 0.000000 40.110000 0.600000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.250000 0.000000 34.390000 0.600000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.530000 0.000000 28.670000 0.600000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.810000 0.000000 22.950000 0.600000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090000 0.000000 17.230000 0.600000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 11.370000 0.000000 11.510000 0.600000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.210000 0.000000 566.350000 0.600000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.490000 0.000000 560.630000 0.600000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.770000 0.000000 554.910000 0.600000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.050000 0.000000 549.190000 0.600000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 543.330000 0.000000 543.470000 0.600000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 537.610000 0.000000 537.750000 0.600000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.890000 0.000000 532.030000 0.600000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.170000 0.000000 526.310000 0.600000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.450000 0.000000 520.590000 0.600000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.730000 0.000000 514.870000 0.600000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.010000 0.000000 509.150000 0.600000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.290000 0.000000 503.430000 0.600000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.570000 0.000000 497.710000 0.600000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.850000 0.000000 491.990000 0.600000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.130000 0.000000 486.270000 0.600000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.410000 0.000000 480.550000 0.600000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.690000 0.000000 474.830000 0.600000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.970000 0.000000 469.110000 0.600000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.250000 0.000000 463.390000 0.600000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.530000 0.000000 457.670000 0.600000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.810000 0.000000 451.950000 0.600000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.090000 0.000000 446.230000 0.600000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 440.370000 0.000000 440.510000 0.600000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.650000 0.000000 434.790000 0.600000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.930000 0.000000 429.070000 0.600000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.210000 0.000000 423.350000 0.600000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 417.490000 0.000000 417.630000 0.600000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 411.770000 0.000000 411.910000 0.600000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.050000 0.000000 406.190000 0.600000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.330000 0.000000 400.470000 0.600000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.610000 0.000000 394.750000 0.600000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 388.890000 0.000000 389.030000 0.600000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1332.690000 0.000000 1332.830000 0.600000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1326.970000 0.000000 1327.110000 0.600000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1321.250000 0.000000 1321.390000 0.600000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1315.530000 0.000000 1315.670000 0.600000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1309.810000 0.000000 1309.950000 0.600000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1304.090000 0.000000 1304.230000 0.600000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1298.370000 0.000000 1298.510000 0.600000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1292.650000 0.000000 1292.790000 0.600000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1286.930000 0.000000 1287.070000 0.600000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1281.210000 0.000000 1281.350000 0.600000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1275.490000 0.000000 1275.630000 0.600000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1269.770000 0.000000 1269.910000 0.600000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1264.050000 0.000000 1264.190000 0.600000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1258.330000 0.000000 1258.470000 0.600000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1252.610000 0.000000 1252.750000 0.600000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1246.890000 0.000000 1247.030000 0.600000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1241.170000 0.000000 1241.310000 0.600000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1235.450000 0.000000 1235.590000 0.600000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1229.730000 0.000000 1229.870000 0.600000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1224.010000 0.000000 1224.150000 0.600000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1218.290000 0.000000 1218.430000 0.600000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1212.570000 0.000000 1212.710000 0.600000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1206.850000 0.000000 1206.990000 0.600000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1201.130000 0.000000 1201.270000 0.600000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1195.410000 0.000000 1195.550000 0.600000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1189.690000 0.000000 1189.830000 0.600000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1183.970000 0.000000 1184.110000 0.600000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1178.250000 0.000000 1178.390000 0.600000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1172.530000 0.000000 1172.670000 0.600000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1166.810000 0.000000 1166.950000 0.600000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1161.090000 0.000000 1161.230000 0.600000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1155.370000 0.000000 1155.510000 0.600000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1149.650000 0.000000 1149.790000 0.600000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1143.930000 0.000000 1144.070000 0.600000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1138.210000 0.000000 1138.350000 0.600000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1132.490000 0.000000 1132.630000 0.600000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1126.770000 0.000000 1126.910000 0.600000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1121.050000 0.000000 1121.190000 0.600000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1115.330000 0.000000 1115.470000 0.600000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1109.610000 0.000000 1109.750000 0.600000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1103.890000 0.000000 1104.030000 0.600000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1098.170000 0.000000 1098.310000 0.600000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1092.450000 0.000000 1092.590000 0.600000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1086.730000 0.000000 1086.870000 0.600000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1081.010000 0.000000 1081.150000 0.600000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1075.290000 0.000000 1075.430000 0.600000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.570000 0.000000 1069.710000 0.600000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.850000 0.000000 1063.990000 0.600000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1058.130000 0.000000 1058.270000 0.600000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1052.410000 0.000000 1052.550000 0.600000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1046.690000 0.000000 1046.830000 0.600000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1040.970000 0.000000 1041.110000 0.600000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.250000 0.000000 1035.390000 0.600000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1029.530000 0.000000 1029.670000 0.600000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1023.810000 0.000000 1023.950000 0.600000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1018.090000 0.000000 1018.230000 0.600000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1012.370000 0.000000 1012.510000 0.600000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1006.650000 0.000000 1006.790000 0.600000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.930000 0.000000 1001.070000 0.600000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 995.210000 0.000000 995.350000 0.600000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 989.490000 0.000000 989.630000 0.600000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 983.770000 0.000000 983.910000 0.600000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 978.050000 0.000000 978.190000 0.600000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.330000 0.000000 972.470000 0.600000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.610000 0.000000 966.750000 0.600000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.890000 0.000000 961.030000 0.600000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 955.170000 0.000000 955.310000 0.600000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 949.450000 0.000000 949.590000 0.600000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 943.730000 0.000000 943.870000 0.600000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.010000 0.000000 938.150000 0.600000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.290000 0.000000 932.430000 0.600000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 926.570000 0.000000 926.710000 0.600000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 920.850000 0.000000 920.990000 0.600000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 915.130000 0.000000 915.270000 0.600000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 909.410000 0.000000 909.550000 0.600000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 903.690000 0.000000 903.830000 0.600000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.970000 0.000000 898.110000 0.600000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 892.250000 0.000000 892.390000 0.600000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 886.530000 0.000000 886.670000 0.600000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 880.810000 0.000000 880.950000 0.600000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 875.090000 0.000000 875.230000 0.600000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.370000 0.000000 869.510000 0.600000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.650000 0.000000 863.790000 0.600000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 857.930000 0.000000 858.070000 0.600000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 852.210000 0.000000 852.350000 0.600000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 846.490000 0.000000 846.630000 0.600000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 840.770000 0.000000 840.910000 0.600000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.050000 0.000000 835.190000 0.600000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 829.330000 0.000000 829.470000 0.600000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 823.610000 0.000000 823.750000 0.600000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 817.890000 0.000000 818.030000 0.600000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 812.170000 0.000000 812.310000 0.600000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 806.450000 0.000000 806.590000 0.600000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.730000 0.000000 800.870000 0.600000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 795.010000 0.000000 795.150000 0.600000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 789.290000 0.000000 789.430000 0.600000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 783.570000 0.000000 783.710000 0.600000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 777.850000 0.000000 777.990000 0.600000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 772.130000 0.000000 772.270000 0.600000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.410000 0.000000 766.550000 0.600000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.690000 0.000000 760.830000 0.600000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 754.970000 0.000000 755.110000 0.600000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 749.250000 0.000000 749.390000 0.600000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 743.530000 0.000000 743.670000 0.600000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 737.810000 0.000000 737.950000 0.600000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.090000 0.000000 732.230000 0.600000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 726.370000 0.000000 726.510000 0.600000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 720.650000 0.000000 720.790000 0.600000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 714.930000 0.000000 715.070000 0.600000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 709.210000 0.000000 709.350000 0.600000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.490000 0.000000 703.630000 0.600000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.770000 0.000000 697.910000 0.600000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 692.050000 0.000000 692.190000 0.600000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 686.330000 0.000000 686.470000 0.600000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 680.610000 0.000000 680.750000 0.600000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 674.890000 0.000000 675.030000 0.600000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.170000 0.000000 669.310000 0.600000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.450000 0.000000 663.590000 0.600000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 657.730000 0.000000 657.870000 0.600000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 652.010000 0.000000 652.150000 0.600000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 646.290000 0.000000 646.430000 0.600000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 640.570000 0.000000 640.710000 0.600000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.850000 0.000000 634.990000 0.600000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.130000 0.000000 629.270000 0.600000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 623.410000 0.000000 623.550000 0.600000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.690000 0.000000 617.830000 0.600000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.970000 0.000000 612.110000 0.600000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.250000 0.000000 606.390000 0.600000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2064.850000 0.000000 2064.990000 0.600000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2059.130000 0.000000 2059.270000 0.600000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2053.410000 0.000000 2053.550000 0.600000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2047.690000 0.000000 2047.830000 0.600000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2041.970000 0.000000 2042.110000 0.600000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2036.250000 0.000000 2036.390000 0.600000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2030.530000 0.000000 2030.670000 0.600000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2024.810000 0.000000 2024.950000 0.600000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2019.090000 0.000000 2019.230000 0.600000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2013.370000 0.000000 2013.510000 0.600000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2007.650000 0.000000 2007.790000 0.600000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2001.930000 0.000000 2002.070000 0.600000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1996.210000 0.000000 1996.350000 0.600000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1990.490000 0.000000 1990.630000 0.600000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1984.770000 0.000000 1984.910000 0.600000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1979.050000 0.000000 1979.190000 0.600000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1973.330000 0.000000 1973.470000 0.600000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1967.610000 0.000000 1967.750000 0.600000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1961.890000 0.000000 1962.030000 0.600000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1956.170000 0.000000 1956.310000 0.600000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1950.450000 0.000000 1950.590000 0.600000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1944.730000 0.000000 1944.870000 0.600000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1939.010000 0.000000 1939.150000 0.600000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1933.290000 0.000000 1933.430000 0.600000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1927.570000 0.000000 1927.710000 0.600000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1921.850000 0.000000 1921.990000 0.600000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1916.130000 0.000000 1916.270000 0.600000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1910.410000 0.000000 1910.550000 0.600000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1904.690000 0.000000 1904.830000 0.600000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1898.970000 0.000000 1899.110000 0.600000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1893.250000 0.000000 1893.390000 0.600000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1887.530000 0.000000 1887.670000 0.600000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1881.810000 0.000000 1881.950000 0.600000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1876.090000 0.000000 1876.230000 0.600000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1870.370000 0.000000 1870.510000 0.600000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1864.650000 0.000000 1864.790000 0.600000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1858.930000 0.000000 1859.070000 0.600000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1853.210000 0.000000 1853.350000 0.600000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1847.490000 0.000000 1847.630000 0.600000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1841.770000 0.000000 1841.910000 0.600000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1836.050000 0.000000 1836.190000 0.600000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1830.330000 0.000000 1830.470000 0.600000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1824.610000 0.000000 1824.750000 0.600000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1818.890000 0.000000 1819.030000 0.600000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1813.170000 0.000000 1813.310000 0.600000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1807.450000 0.000000 1807.590000 0.600000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1801.730000 0.000000 1801.870000 0.600000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1796.010000 0.000000 1796.150000 0.600000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1790.290000 0.000000 1790.430000 0.600000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1784.570000 0.000000 1784.710000 0.600000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1778.850000 0.000000 1778.990000 0.600000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1773.130000 0.000000 1773.270000 0.600000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1767.410000 0.000000 1767.550000 0.600000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1761.690000 0.000000 1761.830000 0.600000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1755.970000 0.000000 1756.110000 0.600000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1750.250000 0.000000 1750.390000 0.600000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1744.530000 0.000000 1744.670000 0.600000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1738.810000 0.000000 1738.950000 0.600000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1733.090000 0.000000 1733.230000 0.600000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1727.370000 0.000000 1727.510000 0.600000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1721.650000 0.000000 1721.790000 0.600000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1715.930000 0.000000 1716.070000 0.600000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1710.210000 0.000000 1710.350000 0.600000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1704.490000 0.000000 1704.630000 0.600000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1698.770000 0.000000 1698.910000 0.600000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1693.050000 0.000000 1693.190000 0.600000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1687.330000 0.000000 1687.470000 0.600000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1681.610000 0.000000 1681.750000 0.600000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1675.890000 0.000000 1676.030000 0.600000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1670.170000 0.000000 1670.310000 0.600000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1664.450000 0.000000 1664.590000 0.600000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1658.730000 0.000000 1658.870000 0.600000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1653.010000 0.000000 1653.150000 0.600000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1647.290000 0.000000 1647.430000 0.600000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1641.570000 0.000000 1641.710000 0.600000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1635.850000 0.000000 1635.990000 0.600000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1630.130000 0.000000 1630.270000 0.600000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1624.410000 0.000000 1624.550000 0.600000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1618.690000 0.000000 1618.830000 0.600000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1612.970000 0.000000 1613.110000 0.600000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1607.250000 0.000000 1607.390000 0.600000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1601.530000 0.000000 1601.670000 0.600000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1595.810000 0.000000 1595.950000 0.600000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1590.090000 0.000000 1590.230000 0.600000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1584.370000 0.000000 1584.510000 0.600000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1578.650000 0.000000 1578.790000 0.600000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1572.930000 0.000000 1573.070000 0.600000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1567.210000 0.000000 1567.350000 0.600000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1561.490000 0.000000 1561.630000 0.600000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1555.770000 0.000000 1555.910000 0.600000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1550.050000 0.000000 1550.190000 0.600000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1544.330000 0.000000 1544.470000 0.600000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1538.610000 0.000000 1538.750000 0.600000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1532.890000 0.000000 1533.030000 0.600000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1527.170000 0.000000 1527.310000 0.600000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1521.450000 0.000000 1521.590000 0.600000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1515.730000 0.000000 1515.870000 0.600000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1510.010000 0.000000 1510.150000 0.600000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1504.290000 0.000000 1504.430000 0.600000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1498.570000 0.000000 1498.710000 0.600000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1492.850000 0.000000 1492.990000 0.600000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1487.130000 0.000000 1487.270000 0.600000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1481.410000 0.000000 1481.550000 0.600000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1475.690000 0.000000 1475.830000 0.600000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1469.970000 0.000000 1470.110000 0.600000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1464.250000 0.000000 1464.390000 0.600000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1458.530000 0.000000 1458.670000 0.600000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1452.810000 0.000000 1452.950000 0.600000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1447.090000 0.000000 1447.230000 0.600000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1441.370000 0.000000 1441.510000 0.600000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1435.650000 0.000000 1435.790000 0.600000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1429.930000 0.000000 1430.070000 0.600000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1424.210000 0.000000 1424.350000 0.600000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.490000 0.000000 1418.630000 0.600000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1412.770000 0.000000 1412.910000 0.600000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1407.050000 0.000000 1407.190000 0.600000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1401.330000 0.000000 1401.470000 0.600000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1395.610000 0.000000 1395.750000 0.600000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1389.890000 0.000000 1390.030000 0.600000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1384.170000 0.000000 1384.310000 0.600000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1378.450000 0.000000 1378.590000 0.600000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1372.730000 0.000000 1372.870000 0.600000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1367.010000 0.000000 1367.150000 0.600000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1361.290000 0.000000 1361.430000 0.600000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1355.570000 0.000000 1355.710000 0.600000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1349.850000 0.000000 1349.990000 0.600000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1344.130000 0.000000 1344.270000 0.600000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.410000 0.000000 1338.550000 0.600000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2797.010000 0.000000 2797.150000 0.600000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2791.290000 0.000000 2791.430000 0.600000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2785.570000 0.000000 2785.710000 0.600000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2779.850000 0.000000 2779.990000 0.600000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2774.130000 0.000000 2774.270000 0.600000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2768.410000 0.000000 2768.550000 0.600000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2762.690000 0.000000 2762.830000 0.600000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2756.970000 0.000000 2757.110000 0.600000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2751.250000 0.000000 2751.390000 0.600000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2745.530000 0.000000 2745.670000 0.600000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2739.810000 0.000000 2739.950000 0.600000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2734.090000 0.000000 2734.230000 0.600000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2728.370000 0.000000 2728.510000 0.600000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2722.650000 0.000000 2722.790000 0.600000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2716.930000 0.000000 2717.070000 0.600000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2711.210000 0.000000 2711.350000 0.600000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2705.490000 0.000000 2705.630000 0.600000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2699.770000 0.000000 2699.910000 0.600000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2694.050000 0.000000 2694.190000 0.600000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2688.330000 0.000000 2688.470000 0.600000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2682.610000 0.000000 2682.750000 0.600000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2676.890000 0.000000 2677.030000 0.600000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2671.170000 0.000000 2671.310000 0.600000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2665.450000 0.000000 2665.590000 0.600000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2659.730000 0.000000 2659.870000 0.600000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2654.010000 0.000000 2654.150000 0.600000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2648.290000 0.000000 2648.430000 0.600000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2642.570000 0.000000 2642.710000 0.600000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2636.850000 0.000000 2636.990000 0.600000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2631.130000 0.000000 2631.270000 0.600000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2625.410000 0.000000 2625.550000 0.600000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.690000 0.000000 2619.830000 0.600000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2613.970000 0.000000 2614.110000 0.600000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2608.250000 0.000000 2608.390000 0.600000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2602.530000 0.000000 2602.670000 0.600000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2596.810000 0.000000 2596.950000 0.600000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2591.090000 0.000000 2591.230000 0.600000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2585.370000 0.000000 2585.510000 0.600000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2579.650000 0.000000 2579.790000 0.600000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2573.930000 0.000000 2574.070000 0.600000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2568.210000 0.000000 2568.350000 0.600000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2562.490000 0.000000 2562.630000 0.600000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2556.770000 0.000000 2556.910000 0.600000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2551.050000 0.000000 2551.190000 0.600000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2545.330000 0.000000 2545.470000 0.600000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2539.610000 0.000000 2539.750000 0.600000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2533.890000 0.000000 2534.030000 0.600000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2528.170000 0.000000 2528.310000 0.600000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2522.450000 0.000000 2522.590000 0.600000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2516.730000 0.000000 2516.870000 0.600000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2511.010000 0.000000 2511.150000 0.600000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2505.290000 0.000000 2505.430000 0.600000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2499.570000 0.000000 2499.710000 0.600000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2493.850000 0.000000 2493.990000 0.600000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2488.130000 0.000000 2488.270000 0.600000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2482.410000 0.000000 2482.550000 0.600000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2476.690000 0.000000 2476.830000 0.600000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2470.970000 0.000000 2471.110000 0.600000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2465.250000 0.000000 2465.390000 0.600000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2459.530000 0.000000 2459.670000 0.600000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2453.810000 0.000000 2453.950000 0.600000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2448.090000 0.000000 2448.230000 0.600000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2442.370000 0.000000 2442.510000 0.600000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2436.650000 0.000000 2436.790000 0.600000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2430.930000 0.000000 2431.070000 0.600000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2425.210000 0.000000 2425.350000 0.600000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2419.490000 0.000000 2419.630000 0.600000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2413.770000 0.000000 2413.910000 0.600000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2408.050000 0.000000 2408.190000 0.600000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2402.330000 0.000000 2402.470000 0.600000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2396.610000 0.000000 2396.750000 0.600000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2390.890000 0.000000 2391.030000 0.600000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2385.170000 0.000000 2385.310000 0.600000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2379.450000 0.000000 2379.590000 0.600000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2373.730000 0.000000 2373.870000 0.600000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2368.010000 0.000000 2368.150000 0.600000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2362.290000 0.000000 2362.430000 0.600000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2356.570000 0.000000 2356.710000 0.600000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2350.850000 0.000000 2350.990000 0.600000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2345.130000 0.000000 2345.270000 0.600000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2339.410000 0.000000 2339.550000 0.600000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2333.690000 0.000000 2333.830000 0.600000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2327.970000 0.000000 2328.110000 0.600000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2322.250000 0.000000 2322.390000 0.600000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2316.530000 0.000000 2316.670000 0.600000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2310.810000 0.000000 2310.950000 0.600000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2305.090000 0.000000 2305.230000 0.600000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2299.370000 0.000000 2299.510000 0.600000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2293.650000 0.000000 2293.790000 0.600000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2287.930000 0.000000 2288.070000 0.600000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2282.210000 0.000000 2282.350000 0.600000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2276.490000 0.000000 2276.630000 0.600000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2270.770000 0.000000 2270.910000 0.600000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2265.050000 0.000000 2265.190000 0.600000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2259.330000 0.000000 2259.470000 0.600000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2253.610000 0.000000 2253.750000 0.600000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2247.890000 0.000000 2248.030000 0.600000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2242.170000 0.000000 2242.310000 0.600000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2236.450000 0.000000 2236.590000 0.600000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2230.730000 0.000000 2230.870000 0.600000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2225.010000 0.000000 2225.150000 0.600000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2219.290000 0.000000 2219.430000 0.600000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2213.570000 0.000000 2213.710000 0.600000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2207.850000 0.000000 2207.990000 0.600000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2202.130000 0.000000 2202.270000 0.600000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2196.410000 0.000000 2196.550000 0.600000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2190.690000 0.000000 2190.830000 0.600000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2184.970000 0.000000 2185.110000 0.600000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2179.250000 0.000000 2179.390000 0.600000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2173.530000 0.000000 2173.670000 0.600000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2167.810000 0.000000 2167.950000 0.600000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2162.090000 0.000000 2162.230000 0.600000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2156.370000 0.000000 2156.510000 0.600000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2150.650000 0.000000 2150.790000 0.600000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2144.930000 0.000000 2145.070000 0.600000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2139.210000 0.000000 2139.350000 0.600000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2133.490000 0.000000 2133.630000 0.600000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2127.770000 0.000000 2127.910000 0.600000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2122.050000 0.000000 2122.190000 0.600000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2116.330000 0.000000 2116.470000 0.600000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2110.610000 0.000000 2110.750000 0.600000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2104.890000 0.000000 2105.030000 0.600000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2099.170000 0.000000 2099.310000 0.600000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2093.450000 0.000000 2093.590000 0.600000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2087.730000 0.000000 2087.870000 0.600000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2082.010000 0.000000 2082.150000 0.600000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2076.290000 0.000000 2076.430000 0.600000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2070.570000 0.000000 2070.710000 0.600000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 121.480000 0.600000 121.620000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 303.720000 0.600000 303.860000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 485.960000 0.600000 486.100000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 729.060000 0.600000 729.200000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 972.160000 0.600000 972.300000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1215.260000 0.600000 1215.400000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1458.020000 0.600000 1458.160000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1701.120000 0.600000 1701.260000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1944.220000 0.600000 1944.360000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2186.980000 0.600000 2187.120000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2430.080000 0.600000 2430.220000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2673.180000 0.600000 2673.320000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2915.940000 0.600000 2916.080000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3159.040000 0.600000 3159.180000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.085000 3219.200000 161.225000 3219.800000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.400000 3219.200000 483.540000 3219.800000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 805.710000 3219.200000 805.850000 3219.800000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1128.020000 3219.200000 1128.160000 3219.800000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1450.335000 3219.200000 1450.475000 3219.800000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1772.645000 3219.200000 1772.785000 3219.800000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2094.960000 3219.200000 2095.100000 3219.800000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2417.270000 3219.200000 2417.410000 3219.800000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2739.580000 3219.200000 2739.720000 3219.800000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 3095.800000 2820.260000 3095.940000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2847.940000 2820.260000 2848.080000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2600.420000 2820.260000 2600.560000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2352.560000 2820.260000 2352.700000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2105.040000 2820.260000 2105.180000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1857.180000 2820.260000 1857.320000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1609.660000 2820.260000 1609.800000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1362.140000 2820.260000 1362.280000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1114.280000 2820.260000 1114.420000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 928.640000 2820.260000 928.780000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 742.660000 2820.260000 742.800000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 557.020000 2820.260000 557.160000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 371.380000 2820.260000 371.520000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 185.400000 2820.260000 185.540000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1.800000 2820.260000 1.940000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 60.960000 0.600000 61.100000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 243.200000 0.600000 243.340000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 425.440000 0.600000 425.580000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 668.200000 0.600000 668.340000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 911.300000 0.600000 911.440000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1154.400000 0.600000 1154.540000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1397.500000 0.600000 1397.640000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1640.260000 0.600000 1640.400000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1883.360000 0.600000 1883.500000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2126.460000 0.600000 2126.600000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2369.220000 0.600000 2369.360000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2612.320000 0.600000 2612.460000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2855.420000 0.600000 2855.560000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3098.180000 0.600000 3098.320000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 80.510000 3219.200000 80.650000 3219.800000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.820000 3219.200000 402.960000 3219.800000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.130000 3219.200000 725.270000 3219.800000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1047.445000 3219.200000 1047.585000 3219.800000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1369.755000 3219.200000 1369.895000 3219.800000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1692.070000 3219.200000 1692.210000 3219.800000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2014.380000 3219.200000 2014.520000 3219.800000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2336.690000 3219.200000 2336.830000 3219.800000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2659.005000 3219.200000 2659.145000 3219.800000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 3157.680000 2820.260000 3157.820000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2909.820000 2820.260000 2909.960000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2662.300000 2820.260000 2662.440000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2414.440000 2820.260000 2414.580000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2166.920000 2820.260000 2167.060000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1919.400000 2820.260000 1919.540000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1671.540000 2820.260000 1671.680000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1424.020000 2820.260000 1424.160000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1176.160000 2820.260000 1176.300000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 990.520000 2820.260000 990.660000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 804.540000 2820.260000 804.680000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 618.900000 2820.260000 619.040000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 433.260000 2820.260000 433.400000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 247.280000 2820.260000 247.420000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 61.640000 2820.260000 61.780000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2.140000 0.600000 2.280000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 182.340000 0.600000 182.480000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 364.580000 0.600000 364.720000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 607.680000 0.600000 607.820000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 850.440000 0.600000 850.580000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1093.540000 0.600000 1093.680000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1336.640000 0.600000 1336.780000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1579.740000 0.600000 1579.880000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1822.500000 0.600000 1822.640000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2065.600000 0.600000 2065.740000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2308.700000 0.600000 2308.840000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2551.460000 0.600000 2551.600000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2794.560000 0.600000 2794.700000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3037.660000 0.600000 3037.800000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.080000 3219.200000 1.220000 3219.800000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 322.240000 3219.200000 322.380000 3219.800000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 644.555000 3219.200000 644.695000 3219.800000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.865000 3219.200000 967.005000 3219.800000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1289.180000 3219.200000 1289.320000 3219.800000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1611.490000 3219.200000 1611.630000 3219.800000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1933.800000 3219.200000 1933.940000 3219.800000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2256.115000 3219.200000 2256.255000 3219.800000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2578.425000 3219.200000 2578.565000 3219.800000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 3214.800000 2820.260000 3214.940000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2972.040000 2820.260000 2972.180000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2724.180000 2820.260000 2724.320000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2476.660000 2820.260000 2476.800000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2228.800000 2820.260000 2228.940000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1981.280000 2820.260000 1981.420000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1733.420000 2820.260000 1733.560000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1485.900000 2820.260000 1486.040000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1238.040000 2820.260000 1238.180000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1052.400000 2820.260000 1052.540000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 866.760000 2820.260000 866.900000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 680.780000 2820.260000 680.920000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 495.140000 2820.260000 495.280000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 309.500000 2820.260000 309.640000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 123.520000 2820.260000 123.660000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 546.820000 0.600000 546.960000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 789.920000 0.600000 790.060000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1032.680000 0.600000 1032.820000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1275.780000 0.600000 1275.920000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1518.880000 0.600000 1519.020000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1761.980000 0.600000 1762.120000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2004.740000 0.600000 2004.880000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2247.840000 0.600000 2247.980000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2490.940000 0.600000 2491.080000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2733.700000 0.600000 2733.840000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2976.800000 0.600000 2976.940000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3215.140000 0.600000 3215.280000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 241.665000 3219.200000 241.805000 3219.800000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 563.975000 3219.200000 564.115000 3219.800000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 886.290000 3219.200000 886.430000 3219.800000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1208.600000 3219.200000 1208.740000 3219.800000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1530.910000 3219.200000 1531.050000 3219.800000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1853.225000 3219.200000 1853.365000 3219.800000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2175.535000 3219.200000 2175.675000 3219.800000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2497.850000 3219.200000 2497.990000 3219.800000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2815.360000 3219.200000 2815.500000 3219.800000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 3033.920000 2820.260000 3034.060000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2786.060000 2820.260000 2786.200000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2538.540000 2820.260000 2538.680000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2290.680000 2820.260000 2290.820000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 2043.160000 2820.260000 2043.300000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1795.300000 2820.260000 1795.440000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1547.780000 2820.260000 1547.920000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.660000 1299.920000 2820.260000 1300.060000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2802.730000 0.000000 2802.870000 0.600000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2819.890000 0.000000 2820.030000 0.600000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2814.170000 0.000000 2814.310000 0.600000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2808.450000 0.000000 2808.590000 0.600000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.160000 1730.487000 4.160000 1742.530000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2005.560000 2696.355000 2007.300000 3091.135000 ;
      LAYER met4 ;
        RECT 1530.240000 2696.355000 1531.980000 3091.135000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1324.945000 2709.480000 1326.685000 3104.260000 ;
      LAYER met4 ;
        RECT 849.625000 2709.480000 851.365000 3104.260000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2649.535000 2700.010000 2651.275000 3094.790000 ;
      LAYER met4 ;
        RECT 2174.215000 2700.010000 2175.955000 3094.790000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 704.015000 2715.950000 705.755000 3110.730000 ;
      LAYER met4 ;
        RECT 228.695000 2715.950000 230.435000 3110.730000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2690.935000 75.330000 2692.675000 470.110000 ;
      LAYER met4 ;
        RECT 2215.615000 75.330000 2217.355000 470.110000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2081.880000 82.810000 2083.620000 477.590000 ;
      LAYER met4 ;
        RECT 1606.560000 82.810000 1608.300000 477.590000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 367.970000 87.900000 369.710000 482.680000 ;
      LAYER met4 ;
        RECT 843.290000 87.900000 845.030000 482.680000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1017.520000 93.075000 1019.260000 487.855000 ;
      LAYER met4 ;
        RECT 1492.840000 93.075000 1494.580000 487.855000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.960000 1716.405000 7.960000 1731.830000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1533.640000 2699.755000 1535.380000 3087.735000 ;
      LAYER met4 ;
        RECT 2002.160000 2699.755000 2003.900000 3087.735000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 853.025000 2712.880000 854.765000 3100.860000 ;
      LAYER met4 ;
        RECT 1321.545000 2712.880000 1323.285000 3100.860000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2177.615000 2703.410000 2179.355000 3091.390000 ;
      LAYER met4 ;
        RECT 2646.135000 2703.410000 2647.875000 3091.390000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 232.095000 2719.350000 233.835000 3107.330000 ;
      LAYER met4 ;
        RECT 700.615000 2719.350000 702.355000 3107.330000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2219.015000 78.730000 2220.755000 466.710000 ;
      LAYER met4 ;
        RECT 2687.535000 78.730000 2689.275000 466.710000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1609.960000 86.210000 1611.700000 474.190000 ;
      LAYER met4 ;
        RECT 2078.480000 86.210000 2080.220000 474.190000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 839.890000 91.300000 841.630000 479.280000 ;
      LAYER met4 ;
        RECT 371.370000 91.300000 373.110000 479.280000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1489.440000 96.475000 1491.180000 484.455000 ;
      LAYER met4 ;
        RECT 1020.920000 96.475000 1022.660000 484.455000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2820.260000 3219.800000 ;
    LAYER met1 ;
      RECT 2815.640000 3219.060000 2820.260000 3219.800000 ;
      RECT 2739.860000 3219.060000 2815.220000 3219.800000 ;
      RECT 2659.285000 3219.060000 2739.440000 3219.800000 ;
      RECT 2578.705000 3219.060000 2658.865000 3219.800000 ;
      RECT 2498.130000 3219.060000 2578.285000 3219.800000 ;
      RECT 2417.550000 3219.060000 2497.710000 3219.800000 ;
      RECT 2336.970000 3219.060000 2417.130000 3219.800000 ;
      RECT 2256.395000 3219.060000 2336.550000 3219.800000 ;
      RECT 2175.815000 3219.060000 2255.975000 3219.800000 ;
      RECT 2095.240000 3219.060000 2175.395000 3219.800000 ;
      RECT 2014.660000 3219.060000 2094.820000 3219.800000 ;
      RECT 1934.080000 3219.060000 2014.240000 3219.800000 ;
      RECT 1853.505000 3219.060000 1933.660000 3219.800000 ;
      RECT 1772.925000 3219.060000 1853.085000 3219.800000 ;
      RECT 1692.350000 3219.060000 1772.505000 3219.800000 ;
      RECT 1611.770000 3219.060000 1691.930000 3219.800000 ;
      RECT 1531.190000 3219.060000 1611.350000 3219.800000 ;
      RECT 1450.615000 3219.060000 1530.770000 3219.800000 ;
      RECT 1370.035000 3219.060000 1450.195000 3219.800000 ;
      RECT 1289.460000 3219.060000 1369.615000 3219.800000 ;
      RECT 1208.880000 3219.060000 1289.040000 3219.800000 ;
      RECT 1128.300000 3219.060000 1208.460000 3219.800000 ;
      RECT 1047.725000 3219.060000 1127.880000 3219.800000 ;
      RECT 967.145000 3219.060000 1047.305000 3219.800000 ;
      RECT 886.570000 3219.060000 966.725000 3219.800000 ;
      RECT 805.990000 3219.060000 886.150000 3219.800000 ;
      RECT 725.410000 3219.060000 805.570000 3219.800000 ;
      RECT 644.835000 3219.060000 724.990000 3219.800000 ;
      RECT 564.255000 3219.060000 644.415000 3219.800000 ;
      RECT 483.680000 3219.060000 563.835000 3219.800000 ;
      RECT 403.100000 3219.060000 483.260000 3219.800000 ;
      RECT 322.520000 3219.060000 402.680000 3219.800000 ;
      RECT 241.945000 3219.060000 322.100000 3219.800000 ;
      RECT 161.365000 3219.060000 241.525000 3219.800000 ;
      RECT 80.790000 3219.060000 160.945000 3219.800000 ;
      RECT 1.360000 3219.060000 80.370000 3219.800000 ;
      RECT 0.000000 3219.060000 0.940000 3219.800000 ;
      RECT 0.000000 0.740000 2820.260000 3219.060000 ;
      RECT 2820.170000 0.000000 2820.260000 0.740000 ;
      RECT 2814.450000 0.000000 2819.750000 0.740000 ;
      RECT 2808.730000 0.000000 2814.030000 0.740000 ;
      RECT 2803.010000 0.000000 2808.310000 0.740000 ;
      RECT 2797.290000 0.000000 2802.590000 0.740000 ;
      RECT 2791.570000 0.000000 2796.870000 0.740000 ;
      RECT 2785.850000 0.000000 2791.150000 0.740000 ;
      RECT 2780.130000 0.000000 2785.430000 0.740000 ;
      RECT 2774.410000 0.000000 2779.710000 0.740000 ;
      RECT 2768.690000 0.000000 2773.990000 0.740000 ;
      RECT 2762.970000 0.000000 2768.270000 0.740000 ;
      RECT 2757.250000 0.000000 2762.550000 0.740000 ;
      RECT 2751.530000 0.000000 2756.830000 0.740000 ;
      RECT 2745.810000 0.000000 2751.110000 0.740000 ;
      RECT 2740.090000 0.000000 2745.390000 0.740000 ;
      RECT 2734.370000 0.000000 2739.670000 0.740000 ;
      RECT 2728.650000 0.000000 2733.950000 0.740000 ;
      RECT 2722.930000 0.000000 2728.230000 0.740000 ;
      RECT 2717.210000 0.000000 2722.510000 0.740000 ;
      RECT 2711.490000 0.000000 2716.790000 0.740000 ;
      RECT 2705.770000 0.000000 2711.070000 0.740000 ;
      RECT 2700.050000 0.000000 2705.350000 0.740000 ;
      RECT 2694.330000 0.000000 2699.630000 0.740000 ;
      RECT 2688.610000 0.000000 2693.910000 0.740000 ;
      RECT 2682.890000 0.000000 2688.190000 0.740000 ;
      RECT 2677.170000 0.000000 2682.470000 0.740000 ;
      RECT 2671.450000 0.000000 2676.750000 0.740000 ;
      RECT 2665.730000 0.000000 2671.030000 0.740000 ;
      RECT 2660.010000 0.000000 2665.310000 0.740000 ;
      RECT 2654.290000 0.000000 2659.590000 0.740000 ;
      RECT 2648.570000 0.000000 2653.870000 0.740000 ;
      RECT 2642.850000 0.000000 2648.150000 0.740000 ;
      RECT 2637.130000 0.000000 2642.430000 0.740000 ;
      RECT 2631.410000 0.000000 2636.710000 0.740000 ;
      RECT 2625.690000 0.000000 2630.990000 0.740000 ;
      RECT 2619.970000 0.000000 2625.270000 0.740000 ;
      RECT 2614.250000 0.000000 2619.550000 0.740000 ;
      RECT 2608.530000 0.000000 2613.830000 0.740000 ;
      RECT 2602.810000 0.000000 2608.110000 0.740000 ;
      RECT 2597.090000 0.000000 2602.390000 0.740000 ;
      RECT 2591.370000 0.000000 2596.670000 0.740000 ;
      RECT 2585.650000 0.000000 2590.950000 0.740000 ;
      RECT 2579.930000 0.000000 2585.230000 0.740000 ;
      RECT 2574.210000 0.000000 2579.510000 0.740000 ;
      RECT 2568.490000 0.000000 2573.790000 0.740000 ;
      RECT 2562.770000 0.000000 2568.070000 0.740000 ;
      RECT 2557.050000 0.000000 2562.350000 0.740000 ;
      RECT 2551.330000 0.000000 2556.630000 0.740000 ;
      RECT 2545.610000 0.000000 2550.910000 0.740000 ;
      RECT 2539.890000 0.000000 2545.190000 0.740000 ;
      RECT 2534.170000 0.000000 2539.470000 0.740000 ;
      RECT 2528.450000 0.000000 2533.750000 0.740000 ;
      RECT 2522.730000 0.000000 2528.030000 0.740000 ;
      RECT 2517.010000 0.000000 2522.310000 0.740000 ;
      RECT 2511.290000 0.000000 2516.590000 0.740000 ;
      RECT 2505.570000 0.000000 2510.870000 0.740000 ;
      RECT 2499.850000 0.000000 2505.150000 0.740000 ;
      RECT 2494.130000 0.000000 2499.430000 0.740000 ;
      RECT 2488.410000 0.000000 2493.710000 0.740000 ;
      RECT 2482.690000 0.000000 2487.990000 0.740000 ;
      RECT 2476.970000 0.000000 2482.270000 0.740000 ;
      RECT 2471.250000 0.000000 2476.550000 0.740000 ;
      RECT 2465.530000 0.000000 2470.830000 0.740000 ;
      RECT 2459.810000 0.000000 2465.110000 0.740000 ;
      RECT 2454.090000 0.000000 2459.390000 0.740000 ;
      RECT 2448.370000 0.000000 2453.670000 0.740000 ;
      RECT 2442.650000 0.000000 2447.950000 0.740000 ;
      RECT 2436.930000 0.000000 2442.230000 0.740000 ;
      RECT 2431.210000 0.000000 2436.510000 0.740000 ;
      RECT 2425.490000 0.000000 2430.790000 0.740000 ;
      RECT 2419.770000 0.000000 2425.070000 0.740000 ;
      RECT 2414.050000 0.000000 2419.350000 0.740000 ;
      RECT 2408.330000 0.000000 2413.630000 0.740000 ;
      RECT 2402.610000 0.000000 2407.910000 0.740000 ;
      RECT 2396.890000 0.000000 2402.190000 0.740000 ;
      RECT 2391.170000 0.000000 2396.470000 0.740000 ;
      RECT 2385.450000 0.000000 2390.750000 0.740000 ;
      RECT 2379.730000 0.000000 2385.030000 0.740000 ;
      RECT 2374.010000 0.000000 2379.310000 0.740000 ;
      RECT 2368.290000 0.000000 2373.590000 0.740000 ;
      RECT 2362.570000 0.000000 2367.870000 0.740000 ;
      RECT 2356.850000 0.000000 2362.150000 0.740000 ;
      RECT 2351.130000 0.000000 2356.430000 0.740000 ;
      RECT 2345.410000 0.000000 2350.710000 0.740000 ;
      RECT 2339.690000 0.000000 2344.990000 0.740000 ;
      RECT 2333.970000 0.000000 2339.270000 0.740000 ;
      RECT 2328.250000 0.000000 2333.550000 0.740000 ;
      RECT 2322.530000 0.000000 2327.830000 0.740000 ;
      RECT 2316.810000 0.000000 2322.110000 0.740000 ;
      RECT 2311.090000 0.000000 2316.390000 0.740000 ;
      RECT 2305.370000 0.000000 2310.670000 0.740000 ;
      RECT 2299.650000 0.000000 2304.950000 0.740000 ;
      RECT 2293.930000 0.000000 2299.230000 0.740000 ;
      RECT 2288.210000 0.000000 2293.510000 0.740000 ;
      RECT 2282.490000 0.000000 2287.790000 0.740000 ;
      RECT 2276.770000 0.000000 2282.070000 0.740000 ;
      RECT 2271.050000 0.000000 2276.350000 0.740000 ;
      RECT 2265.330000 0.000000 2270.630000 0.740000 ;
      RECT 2259.610000 0.000000 2264.910000 0.740000 ;
      RECT 2253.890000 0.000000 2259.190000 0.740000 ;
      RECT 2248.170000 0.000000 2253.470000 0.740000 ;
      RECT 2242.450000 0.000000 2247.750000 0.740000 ;
      RECT 2236.730000 0.000000 2242.030000 0.740000 ;
      RECT 2231.010000 0.000000 2236.310000 0.740000 ;
      RECT 2225.290000 0.000000 2230.590000 0.740000 ;
      RECT 2219.570000 0.000000 2224.870000 0.740000 ;
      RECT 2213.850000 0.000000 2219.150000 0.740000 ;
      RECT 2208.130000 0.000000 2213.430000 0.740000 ;
      RECT 2202.410000 0.000000 2207.710000 0.740000 ;
      RECT 2196.690000 0.000000 2201.990000 0.740000 ;
      RECT 2190.970000 0.000000 2196.270000 0.740000 ;
      RECT 2185.250000 0.000000 2190.550000 0.740000 ;
      RECT 2179.530000 0.000000 2184.830000 0.740000 ;
      RECT 2173.810000 0.000000 2179.110000 0.740000 ;
      RECT 2168.090000 0.000000 2173.390000 0.740000 ;
      RECT 2162.370000 0.000000 2167.670000 0.740000 ;
      RECT 2156.650000 0.000000 2161.950000 0.740000 ;
      RECT 2150.930000 0.000000 2156.230000 0.740000 ;
      RECT 2145.210000 0.000000 2150.510000 0.740000 ;
      RECT 2139.490000 0.000000 2144.790000 0.740000 ;
      RECT 2133.770000 0.000000 2139.070000 0.740000 ;
      RECT 2128.050000 0.000000 2133.350000 0.740000 ;
      RECT 2122.330000 0.000000 2127.630000 0.740000 ;
      RECT 2116.610000 0.000000 2121.910000 0.740000 ;
      RECT 2110.890000 0.000000 2116.190000 0.740000 ;
      RECT 2105.170000 0.000000 2110.470000 0.740000 ;
      RECT 2099.450000 0.000000 2104.750000 0.740000 ;
      RECT 2093.730000 0.000000 2099.030000 0.740000 ;
      RECT 2088.010000 0.000000 2093.310000 0.740000 ;
      RECT 2082.290000 0.000000 2087.590000 0.740000 ;
      RECT 2076.570000 0.000000 2081.870000 0.740000 ;
      RECT 2070.850000 0.000000 2076.150000 0.740000 ;
      RECT 2065.130000 0.000000 2070.430000 0.740000 ;
      RECT 2059.410000 0.000000 2064.710000 0.740000 ;
      RECT 2053.690000 0.000000 2058.990000 0.740000 ;
      RECT 2047.970000 0.000000 2053.270000 0.740000 ;
      RECT 2042.250000 0.000000 2047.550000 0.740000 ;
      RECT 2036.530000 0.000000 2041.830000 0.740000 ;
      RECT 2030.810000 0.000000 2036.110000 0.740000 ;
      RECT 2025.090000 0.000000 2030.390000 0.740000 ;
      RECT 2019.370000 0.000000 2024.670000 0.740000 ;
      RECT 2013.650000 0.000000 2018.950000 0.740000 ;
      RECT 2007.930000 0.000000 2013.230000 0.740000 ;
      RECT 2002.210000 0.000000 2007.510000 0.740000 ;
      RECT 1996.490000 0.000000 2001.790000 0.740000 ;
      RECT 1990.770000 0.000000 1996.070000 0.740000 ;
      RECT 1985.050000 0.000000 1990.350000 0.740000 ;
      RECT 1979.330000 0.000000 1984.630000 0.740000 ;
      RECT 1973.610000 0.000000 1978.910000 0.740000 ;
      RECT 1967.890000 0.000000 1973.190000 0.740000 ;
      RECT 1962.170000 0.000000 1967.470000 0.740000 ;
      RECT 1956.450000 0.000000 1961.750000 0.740000 ;
      RECT 1950.730000 0.000000 1956.030000 0.740000 ;
      RECT 1945.010000 0.000000 1950.310000 0.740000 ;
      RECT 1939.290000 0.000000 1944.590000 0.740000 ;
      RECT 1933.570000 0.000000 1938.870000 0.740000 ;
      RECT 1927.850000 0.000000 1933.150000 0.740000 ;
      RECT 1922.130000 0.000000 1927.430000 0.740000 ;
      RECT 1916.410000 0.000000 1921.710000 0.740000 ;
      RECT 1910.690000 0.000000 1915.990000 0.740000 ;
      RECT 1904.970000 0.000000 1910.270000 0.740000 ;
      RECT 1899.250000 0.000000 1904.550000 0.740000 ;
      RECT 1893.530000 0.000000 1898.830000 0.740000 ;
      RECT 1887.810000 0.000000 1893.110000 0.740000 ;
      RECT 1882.090000 0.000000 1887.390000 0.740000 ;
      RECT 1876.370000 0.000000 1881.670000 0.740000 ;
      RECT 1870.650000 0.000000 1875.950000 0.740000 ;
      RECT 1864.930000 0.000000 1870.230000 0.740000 ;
      RECT 1859.210000 0.000000 1864.510000 0.740000 ;
      RECT 1853.490000 0.000000 1858.790000 0.740000 ;
      RECT 1847.770000 0.000000 1853.070000 0.740000 ;
      RECT 1842.050000 0.000000 1847.350000 0.740000 ;
      RECT 1836.330000 0.000000 1841.630000 0.740000 ;
      RECT 1830.610000 0.000000 1835.910000 0.740000 ;
      RECT 1824.890000 0.000000 1830.190000 0.740000 ;
      RECT 1819.170000 0.000000 1824.470000 0.740000 ;
      RECT 1813.450000 0.000000 1818.750000 0.740000 ;
      RECT 1807.730000 0.000000 1813.030000 0.740000 ;
      RECT 1802.010000 0.000000 1807.310000 0.740000 ;
      RECT 1796.290000 0.000000 1801.590000 0.740000 ;
      RECT 1790.570000 0.000000 1795.870000 0.740000 ;
      RECT 1784.850000 0.000000 1790.150000 0.740000 ;
      RECT 1779.130000 0.000000 1784.430000 0.740000 ;
      RECT 1773.410000 0.000000 1778.710000 0.740000 ;
      RECT 1767.690000 0.000000 1772.990000 0.740000 ;
      RECT 1761.970000 0.000000 1767.270000 0.740000 ;
      RECT 1756.250000 0.000000 1761.550000 0.740000 ;
      RECT 1750.530000 0.000000 1755.830000 0.740000 ;
      RECT 1744.810000 0.000000 1750.110000 0.740000 ;
      RECT 1739.090000 0.000000 1744.390000 0.740000 ;
      RECT 1733.370000 0.000000 1738.670000 0.740000 ;
      RECT 1727.650000 0.000000 1732.950000 0.740000 ;
      RECT 1721.930000 0.000000 1727.230000 0.740000 ;
      RECT 1716.210000 0.000000 1721.510000 0.740000 ;
      RECT 1710.490000 0.000000 1715.790000 0.740000 ;
      RECT 1704.770000 0.000000 1710.070000 0.740000 ;
      RECT 1699.050000 0.000000 1704.350000 0.740000 ;
      RECT 1693.330000 0.000000 1698.630000 0.740000 ;
      RECT 1687.610000 0.000000 1692.910000 0.740000 ;
      RECT 1681.890000 0.000000 1687.190000 0.740000 ;
      RECT 1676.170000 0.000000 1681.470000 0.740000 ;
      RECT 1670.450000 0.000000 1675.750000 0.740000 ;
      RECT 1664.730000 0.000000 1670.030000 0.740000 ;
      RECT 1659.010000 0.000000 1664.310000 0.740000 ;
      RECT 1653.290000 0.000000 1658.590000 0.740000 ;
      RECT 1647.570000 0.000000 1652.870000 0.740000 ;
      RECT 1641.850000 0.000000 1647.150000 0.740000 ;
      RECT 1636.130000 0.000000 1641.430000 0.740000 ;
      RECT 1630.410000 0.000000 1635.710000 0.740000 ;
      RECT 1624.690000 0.000000 1629.990000 0.740000 ;
      RECT 1618.970000 0.000000 1624.270000 0.740000 ;
      RECT 1613.250000 0.000000 1618.550000 0.740000 ;
      RECT 1607.530000 0.000000 1612.830000 0.740000 ;
      RECT 1601.810000 0.000000 1607.110000 0.740000 ;
      RECT 1596.090000 0.000000 1601.390000 0.740000 ;
      RECT 1590.370000 0.000000 1595.670000 0.740000 ;
      RECT 1584.650000 0.000000 1589.950000 0.740000 ;
      RECT 1578.930000 0.000000 1584.230000 0.740000 ;
      RECT 1573.210000 0.000000 1578.510000 0.740000 ;
      RECT 1567.490000 0.000000 1572.790000 0.740000 ;
      RECT 1561.770000 0.000000 1567.070000 0.740000 ;
      RECT 1556.050000 0.000000 1561.350000 0.740000 ;
      RECT 1550.330000 0.000000 1555.630000 0.740000 ;
      RECT 1544.610000 0.000000 1549.910000 0.740000 ;
      RECT 1538.890000 0.000000 1544.190000 0.740000 ;
      RECT 1533.170000 0.000000 1538.470000 0.740000 ;
      RECT 1527.450000 0.000000 1532.750000 0.740000 ;
      RECT 1521.730000 0.000000 1527.030000 0.740000 ;
      RECT 1516.010000 0.000000 1521.310000 0.740000 ;
      RECT 1510.290000 0.000000 1515.590000 0.740000 ;
      RECT 1504.570000 0.000000 1509.870000 0.740000 ;
      RECT 1498.850000 0.000000 1504.150000 0.740000 ;
      RECT 1493.130000 0.000000 1498.430000 0.740000 ;
      RECT 1487.410000 0.000000 1492.710000 0.740000 ;
      RECT 1481.690000 0.000000 1486.990000 0.740000 ;
      RECT 1475.970000 0.000000 1481.270000 0.740000 ;
      RECT 1470.250000 0.000000 1475.550000 0.740000 ;
      RECT 1464.530000 0.000000 1469.830000 0.740000 ;
      RECT 1458.810000 0.000000 1464.110000 0.740000 ;
      RECT 1453.090000 0.000000 1458.390000 0.740000 ;
      RECT 1447.370000 0.000000 1452.670000 0.740000 ;
      RECT 1441.650000 0.000000 1446.950000 0.740000 ;
      RECT 1435.930000 0.000000 1441.230000 0.740000 ;
      RECT 1430.210000 0.000000 1435.510000 0.740000 ;
      RECT 1424.490000 0.000000 1429.790000 0.740000 ;
      RECT 1418.770000 0.000000 1424.070000 0.740000 ;
      RECT 1413.050000 0.000000 1418.350000 0.740000 ;
      RECT 1407.330000 0.000000 1412.630000 0.740000 ;
      RECT 1401.610000 0.000000 1406.910000 0.740000 ;
      RECT 1395.890000 0.000000 1401.190000 0.740000 ;
      RECT 1390.170000 0.000000 1395.470000 0.740000 ;
      RECT 1384.450000 0.000000 1389.750000 0.740000 ;
      RECT 1378.730000 0.000000 1384.030000 0.740000 ;
      RECT 1373.010000 0.000000 1378.310000 0.740000 ;
      RECT 1367.290000 0.000000 1372.590000 0.740000 ;
      RECT 1361.570000 0.000000 1366.870000 0.740000 ;
      RECT 1355.850000 0.000000 1361.150000 0.740000 ;
      RECT 1350.130000 0.000000 1355.430000 0.740000 ;
      RECT 1344.410000 0.000000 1349.710000 0.740000 ;
      RECT 1338.690000 0.000000 1343.990000 0.740000 ;
      RECT 1332.970000 0.000000 1338.270000 0.740000 ;
      RECT 1327.250000 0.000000 1332.550000 0.740000 ;
      RECT 1321.530000 0.000000 1326.830000 0.740000 ;
      RECT 1315.810000 0.000000 1321.110000 0.740000 ;
      RECT 1310.090000 0.000000 1315.390000 0.740000 ;
      RECT 1304.370000 0.000000 1309.670000 0.740000 ;
      RECT 1298.650000 0.000000 1303.950000 0.740000 ;
      RECT 1292.930000 0.000000 1298.230000 0.740000 ;
      RECT 1287.210000 0.000000 1292.510000 0.740000 ;
      RECT 1281.490000 0.000000 1286.790000 0.740000 ;
      RECT 1275.770000 0.000000 1281.070000 0.740000 ;
      RECT 1270.050000 0.000000 1275.350000 0.740000 ;
      RECT 1264.330000 0.000000 1269.630000 0.740000 ;
      RECT 1258.610000 0.000000 1263.910000 0.740000 ;
      RECT 1252.890000 0.000000 1258.190000 0.740000 ;
      RECT 1247.170000 0.000000 1252.470000 0.740000 ;
      RECT 1241.450000 0.000000 1246.750000 0.740000 ;
      RECT 1235.730000 0.000000 1241.030000 0.740000 ;
      RECT 1230.010000 0.000000 1235.310000 0.740000 ;
      RECT 1224.290000 0.000000 1229.590000 0.740000 ;
      RECT 1218.570000 0.000000 1223.870000 0.740000 ;
      RECT 1212.850000 0.000000 1218.150000 0.740000 ;
      RECT 1207.130000 0.000000 1212.430000 0.740000 ;
      RECT 1201.410000 0.000000 1206.710000 0.740000 ;
      RECT 1195.690000 0.000000 1200.990000 0.740000 ;
      RECT 1189.970000 0.000000 1195.270000 0.740000 ;
      RECT 1184.250000 0.000000 1189.550000 0.740000 ;
      RECT 1178.530000 0.000000 1183.830000 0.740000 ;
      RECT 1172.810000 0.000000 1178.110000 0.740000 ;
      RECT 1167.090000 0.000000 1172.390000 0.740000 ;
      RECT 1161.370000 0.000000 1166.670000 0.740000 ;
      RECT 1155.650000 0.000000 1160.950000 0.740000 ;
      RECT 1149.930000 0.000000 1155.230000 0.740000 ;
      RECT 1144.210000 0.000000 1149.510000 0.740000 ;
      RECT 1138.490000 0.000000 1143.790000 0.740000 ;
      RECT 1132.770000 0.000000 1138.070000 0.740000 ;
      RECT 1127.050000 0.000000 1132.350000 0.740000 ;
      RECT 1121.330000 0.000000 1126.630000 0.740000 ;
      RECT 1115.610000 0.000000 1120.910000 0.740000 ;
      RECT 1109.890000 0.000000 1115.190000 0.740000 ;
      RECT 1104.170000 0.000000 1109.470000 0.740000 ;
      RECT 1098.450000 0.000000 1103.750000 0.740000 ;
      RECT 1092.730000 0.000000 1098.030000 0.740000 ;
      RECT 1087.010000 0.000000 1092.310000 0.740000 ;
      RECT 1081.290000 0.000000 1086.590000 0.740000 ;
      RECT 1075.570000 0.000000 1080.870000 0.740000 ;
      RECT 1069.850000 0.000000 1075.150000 0.740000 ;
      RECT 1064.130000 0.000000 1069.430000 0.740000 ;
      RECT 1058.410000 0.000000 1063.710000 0.740000 ;
      RECT 1052.690000 0.000000 1057.990000 0.740000 ;
      RECT 1046.970000 0.000000 1052.270000 0.740000 ;
      RECT 1041.250000 0.000000 1046.550000 0.740000 ;
      RECT 1035.530000 0.000000 1040.830000 0.740000 ;
      RECT 1029.810000 0.000000 1035.110000 0.740000 ;
      RECT 1024.090000 0.000000 1029.390000 0.740000 ;
      RECT 1018.370000 0.000000 1023.670000 0.740000 ;
      RECT 1012.650000 0.000000 1017.950000 0.740000 ;
      RECT 1006.930000 0.000000 1012.230000 0.740000 ;
      RECT 1001.210000 0.000000 1006.510000 0.740000 ;
      RECT 995.490000 0.000000 1000.790000 0.740000 ;
      RECT 989.770000 0.000000 995.070000 0.740000 ;
      RECT 984.050000 0.000000 989.350000 0.740000 ;
      RECT 978.330000 0.000000 983.630000 0.740000 ;
      RECT 972.610000 0.000000 977.910000 0.740000 ;
      RECT 966.890000 0.000000 972.190000 0.740000 ;
      RECT 961.170000 0.000000 966.470000 0.740000 ;
      RECT 955.450000 0.000000 960.750000 0.740000 ;
      RECT 949.730000 0.000000 955.030000 0.740000 ;
      RECT 944.010000 0.000000 949.310000 0.740000 ;
      RECT 938.290000 0.000000 943.590000 0.740000 ;
      RECT 932.570000 0.000000 937.870000 0.740000 ;
      RECT 926.850000 0.000000 932.150000 0.740000 ;
      RECT 921.130000 0.000000 926.430000 0.740000 ;
      RECT 915.410000 0.000000 920.710000 0.740000 ;
      RECT 909.690000 0.000000 914.990000 0.740000 ;
      RECT 903.970000 0.000000 909.270000 0.740000 ;
      RECT 898.250000 0.000000 903.550000 0.740000 ;
      RECT 892.530000 0.000000 897.830000 0.740000 ;
      RECT 886.810000 0.000000 892.110000 0.740000 ;
      RECT 881.090000 0.000000 886.390000 0.740000 ;
      RECT 875.370000 0.000000 880.670000 0.740000 ;
      RECT 869.650000 0.000000 874.950000 0.740000 ;
      RECT 863.930000 0.000000 869.230000 0.740000 ;
      RECT 858.210000 0.000000 863.510000 0.740000 ;
      RECT 852.490000 0.000000 857.790000 0.740000 ;
      RECT 846.770000 0.000000 852.070000 0.740000 ;
      RECT 841.050000 0.000000 846.350000 0.740000 ;
      RECT 835.330000 0.000000 840.630000 0.740000 ;
      RECT 829.610000 0.000000 834.910000 0.740000 ;
      RECT 823.890000 0.000000 829.190000 0.740000 ;
      RECT 818.170000 0.000000 823.470000 0.740000 ;
      RECT 812.450000 0.000000 817.750000 0.740000 ;
      RECT 806.730000 0.000000 812.030000 0.740000 ;
      RECT 801.010000 0.000000 806.310000 0.740000 ;
      RECT 795.290000 0.000000 800.590000 0.740000 ;
      RECT 789.570000 0.000000 794.870000 0.740000 ;
      RECT 783.850000 0.000000 789.150000 0.740000 ;
      RECT 778.130000 0.000000 783.430000 0.740000 ;
      RECT 772.410000 0.000000 777.710000 0.740000 ;
      RECT 766.690000 0.000000 771.990000 0.740000 ;
      RECT 760.970000 0.000000 766.270000 0.740000 ;
      RECT 755.250000 0.000000 760.550000 0.740000 ;
      RECT 749.530000 0.000000 754.830000 0.740000 ;
      RECT 743.810000 0.000000 749.110000 0.740000 ;
      RECT 738.090000 0.000000 743.390000 0.740000 ;
      RECT 732.370000 0.000000 737.670000 0.740000 ;
      RECT 726.650000 0.000000 731.950000 0.740000 ;
      RECT 720.930000 0.000000 726.230000 0.740000 ;
      RECT 715.210000 0.000000 720.510000 0.740000 ;
      RECT 709.490000 0.000000 714.790000 0.740000 ;
      RECT 703.770000 0.000000 709.070000 0.740000 ;
      RECT 698.050000 0.000000 703.350000 0.740000 ;
      RECT 692.330000 0.000000 697.630000 0.740000 ;
      RECT 686.610000 0.000000 691.910000 0.740000 ;
      RECT 680.890000 0.000000 686.190000 0.740000 ;
      RECT 675.170000 0.000000 680.470000 0.740000 ;
      RECT 669.450000 0.000000 674.750000 0.740000 ;
      RECT 663.730000 0.000000 669.030000 0.740000 ;
      RECT 658.010000 0.000000 663.310000 0.740000 ;
      RECT 652.290000 0.000000 657.590000 0.740000 ;
      RECT 646.570000 0.000000 651.870000 0.740000 ;
      RECT 640.850000 0.000000 646.150000 0.740000 ;
      RECT 635.130000 0.000000 640.430000 0.740000 ;
      RECT 629.410000 0.000000 634.710000 0.740000 ;
      RECT 623.690000 0.000000 628.990000 0.740000 ;
      RECT 617.970000 0.000000 623.270000 0.740000 ;
      RECT 612.250000 0.000000 617.550000 0.740000 ;
      RECT 606.530000 0.000000 611.830000 0.740000 ;
      RECT 600.810000 0.000000 606.110000 0.740000 ;
      RECT 595.090000 0.000000 600.390000 0.740000 ;
      RECT 589.370000 0.000000 594.670000 0.740000 ;
      RECT 583.650000 0.000000 588.950000 0.740000 ;
      RECT 577.930000 0.000000 583.230000 0.740000 ;
      RECT 572.210000 0.000000 577.510000 0.740000 ;
      RECT 566.490000 0.000000 571.790000 0.740000 ;
      RECT 560.770000 0.000000 566.070000 0.740000 ;
      RECT 555.050000 0.000000 560.350000 0.740000 ;
      RECT 549.330000 0.000000 554.630000 0.740000 ;
      RECT 543.610000 0.000000 548.910000 0.740000 ;
      RECT 537.890000 0.000000 543.190000 0.740000 ;
      RECT 532.170000 0.000000 537.470000 0.740000 ;
      RECT 526.450000 0.000000 531.750000 0.740000 ;
      RECT 520.730000 0.000000 526.030000 0.740000 ;
      RECT 515.010000 0.000000 520.310000 0.740000 ;
      RECT 509.290000 0.000000 514.590000 0.740000 ;
      RECT 503.570000 0.000000 508.870000 0.740000 ;
      RECT 497.850000 0.000000 503.150000 0.740000 ;
      RECT 492.130000 0.000000 497.430000 0.740000 ;
      RECT 486.410000 0.000000 491.710000 0.740000 ;
      RECT 480.690000 0.000000 485.990000 0.740000 ;
      RECT 474.970000 0.000000 480.270000 0.740000 ;
      RECT 469.250000 0.000000 474.550000 0.740000 ;
      RECT 463.530000 0.000000 468.830000 0.740000 ;
      RECT 457.810000 0.000000 463.110000 0.740000 ;
      RECT 452.090000 0.000000 457.390000 0.740000 ;
      RECT 446.370000 0.000000 451.670000 0.740000 ;
      RECT 440.650000 0.000000 445.950000 0.740000 ;
      RECT 434.930000 0.000000 440.230000 0.740000 ;
      RECT 429.210000 0.000000 434.510000 0.740000 ;
      RECT 423.490000 0.000000 428.790000 0.740000 ;
      RECT 417.770000 0.000000 423.070000 0.740000 ;
      RECT 412.050000 0.000000 417.350000 0.740000 ;
      RECT 406.330000 0.000000 411.630000 0.740000 ;
      RECT 400.610000 0.000000 405.910000 0.740000 ;
      RECT 394.890000 0.000000 400.190000 0.740000 ;
      RECT 389.170000 0.000000 394.470000 0.740000 ;
      RECT 383.450000 0.000000 388.750000 0.740000 ;
      RECT 377.730000 0.000000 383.030000 0.740000 ;
      RECT 372.010000 0.000000 377.310000 0.740000 ;
      RECT 366.290000 0.000000 371.590000 0.740000 ;
      RECT 360.570000 0.000000 365.870000 0.740000 ;
      RECT 354.850000 0.000000 360.150000 0.740000 ;
      RECT 349.130000 0.000000 354.430000 0.740000 ;
      RECT 343.410000 0.000000 348.710000 0.740000 ;
      RECT 337.690000 0.000000 342.990000 0.740000 ;
      RECT 331.970000 0.000000 337.270000 0.740000 ;
      RECT 326.250000 0.000000 331.550000 0.740000 ;
      RECT 320.530000 0.000000 325.830000 0.740000 ;
      RECT 314.810000 0.000000 320.110000 0.740000 ;
      RECT 309.090000 0.000000 314.390000 0.740000 ;
      RECT 303.370000 0.000000 308.670000 0.740000 ;
      RECT 297.650000 0.000000 302.950000 0.740000 ;
      RECT 291.930000 0.000000 297.230000 0.740000 ;
      RECT 286.210000 0.000000 291.510000 0.740000 ;
      RECT 280.490000 0.000000 285.790000 0.740000 ;
      RECT 274.770000 0.000000 280.070000 0.740000 ;
      RECT 269.050000 0.000000 274.350000 0.740000 ;
      RECT 263.330000 0.000000 268.630000 0.740000 ;
      RECT 257.610000 0.000000 262.910000 0.740000 ;
      RECT 251.890000 0.000000 257.190000 0.740000 ;
      RECT 246.170000 0.000000 251.470000 0.740000 ;
      RECT 240.450000 0.000000 245.750000 0.740000 ;
      RECT 234.730000 0.000000 240.030000 0.740000 ;
      RECT 229.010000 0.000000 234.310000 0.740000 ;
      RECT 223.290000 0.000000 228.590000 0.740000 ;
      RECT 217.570000 0.000000 222.870000 0.740000 ;
      RECT 211.850000 0.000000 217.150000 0.740000 ;
      RECT 206.130000 0.000000 211.430000 0.740000 ;
      RECT 200.410000 0.000000 205.710000 0.740000 ;
      RECT 194.690000 0.000000 199.990000 0.740000 ;
      RECT 188.970000 0.000000 194.270000 0.740000 ;
      RECT 183.250000 0.000000 188.550000 0.740000 ;
      RECT 177.530000 0.000000 182.830000 0.740000 ;
      RECT 171.810000 0.000000 177.110000 0.740000 ;
      RECT 166.090000 0.000000 171.390000 0.740000 ;
      RECT 160.370000 0.000000 165.670000 0.740000 ;
      RECT 154.650000 0.000000 159.950000 0.740000 ;
      RECT 148.930000 0.000000 154.230000 0.740000 ;
      RECT 143.210000 0.000000 148.510000 0.740000 ;
      RECT 137.490000 0.000000 142.790000 0.740000 ;
      RECT 131.770000 0.000000 137.070000 0.740000 ;
      RECT 126.050000 0.000000 131.350000 0.740000 ;
      RECT 120.330000 0.000000 125.630000 0.740000 ;
      RECT 114.610000 0.000000 119.910000 0.740000 ;
      RECT 108.890000 0.000000 114.190000 0.740000 ;
      RECT 103.170000 0.000000 108.470000 0.740000 ;
      RECT 97.450000 0.000000 102.750000 0.740000 ;
      RECT 91.730000 0.000000 97.030000 0.740000 ;
      RECT 86.010000 0.000000 91.310000 0.740000 ;
      RECT 80.290000 0.000000 85.590000 0.740000 ;
      RECT 74.570000 0.000000 79.870000 0.740000 ;
      RECT 68.850000 0.000000 74.150000 0.740000 ;
      RECT 63.130000 0.000000 68.430000 0.740000 ;
      RECT 57.410000 0.000000 62.710000 0.740000 ;
      RECT 51.690000 0.000000 56.990000 0.740000 ;
      RECT 45.970000 0.000000 51.270000 0.740000 ;
      RECT 40.250000 0.000000 45.550000 0.740000 ;
      RECT 34.530000 0.000000 39.830000 0.740000 ;
      RECT 28.810000 0.000000 34.110000 0.740000 ;
      RECT 23.090000 0.000000 28.390000 0.740000 ;
      RECT 17.370000 0.000000 22.670000 0.740000 ;
      RECT 11.650000 0.000000 16.950000 0.740000 ;
      RECT 5.930000 0.000000 11.230000 0.740000 ;
      RECT 1.820000 0.000000 5.510000 0.740000 ;
      RECT 0.000000 0.000000 1.400000 0.740000 ;
    LAYER met2 ;
      RECT 0.000000 3215.420000 2820.260000 3219.800000 ;
      RECT 0.740000 3215.080000 2820.260000 3215.420000 ;
      RECT 0.740000 3215.000000 2819.520000 3215.080000 ;
      RECT 0.000000 3214.660000 2819.520000 3215.000000 ;
      RECT 0.000000 3159.320000 2820.260000 3214.660000 ;
      RECT 0.740000 3158.900000 2820.260000 3159.320000 ;
      RECT 0.000000 3157.960000 2820.260000 3158.900000 ;
      RECT 0.000000 3157.540000 2819.520000 3157.960000 ;
      RECT 0.000000 3098.460000 2820.260000 3157.540000 ;
      RECT 0.740000 3098.040000 2820.260000 3098.460000 ;
      RECT 0.000000 3096.080000 2820.260000 3098.040000 ;
      RECT 0.000000 3095.660000 2819.520000 3096.080000 ;
      RECT 0.000000 3037.940000 2820.260000 3095.660000 ;
      RECT 0.740000 3037.520000 2820.260000 3037.940000 ;
      RECT 0.000000 3034.200000 2820.260000 3037.520000 ;
      RECT 0.000000 3033.780000 2819.520000 3034.200000 ;
      RECT 0.000000 2977.080000 2820.260000 3033.780000 ;
      RECT 0.740000 2976.660000 2820.260000 2977.080000 ;
      RECT 0.000000 2972.320000 2820.260000 2976.660000 ;
      RECT 0.000000 2971.900000 2819.520000 2972.320000 ;
      RECT 0.000000 2916.220000 2820.260000 2971.900000 ;
      RECT 0.740000 2915.800000 2820.260000 2916.220000 ;
      RECT 0.000000 2910.100000 2820.260000 2915.800000 ;
      RECT 0.000000 2909.680000 2819.520000 2910.100000 ;
      RECT 0.000000 2855.700000 2820.260000 2909.680000 ;
      RECT 0.740000 2855.280000 2820.260000 2855.700000 ;
      RECT 0.000000 2848.220000 2820.260000 2855.280000 ;
      RECT 0.000000 2847.800000 2819.520000 2848.220000 ;
      RECT 0.000000 2794.840000 2820.260000 2847.800000 ;
      RECT 0.740000 2794.420000 2820.260000 2794.840000 ;
      RECT 0.000000 2786.340000 2820.260000 2794.420000 ;
      RECT 0.000000 2785.920000 2819.520000 2786.340000 ;
      RECT 0.000000 2733.980000 2820.260000 2785.920000 ;
      RECT 0.740000 2733.560000 2820.260000 2733.980000 ;
      RECT 0.000000 2724.460000 2820.260000 2733.560000 ;
      RECT 0.000000 2724.040000 2819.520000 2724.460000 ;
      RECT 0.000000 2673.460000 2820.260000 2724.040000 ;
      RECT 0.740000 2673.040000 2820.260000 2673.460000 ;
      RECT 0.000000 2662.580000 2820.260000 2673.040000 ;
      RECT 0.000000 2662.160000 2819.520000 2662.580000 ;
      RECT 0.000000 2612.600000 2820.260000 2662.160000 ;
      RECT 0.740000 2612.180000 2820.260000 2612.600000 ;
      RECT 0.000000 2600.700000 2820.260000 2612.180000 ;
      RECT 0.000000 2600.280000 2819.520000 2600.700000 ;
      RECT 0.000000 2551.740000 2820.260000 2600.280000 ;
      RECT 0.740000 2551.320000 2820.260000 2551.740000 ;
      RECT 0.000000 2538.820000 2820.260000 2551.320000 ;
      RECT 0.000000 2538.400000 2819.520000 2538.820000 ;
      RECT 0.000000 2491.220000 2820.260000 2538.400000 ;
      RECT 0.740000 2490.800000 2820.260000 2491.220000 ;
      RECT 0.000000 2476.940000 2820.260000 2490.800000 ;
      RECT 0.000000 2476.520000 2819.520000 2476.940000 ;
      RECT 0.000000 2430.360000 2820.260000 2476.520000 ;
      RECT 0.740000 2429.940000 2820.260000 2430.360000 ;
      RECT 0.000000 2414.720000 2820.260000 2429.940000 ;
      RECT 0.000000 2414.300000 2819.520000 2414.720000 ;
      RECT 0.000000 2369.500000 2820.260000 2414.300000 ;
      RECT 0.740000 2369.080000 2820.260000 2369.500000 ;
      RECT 0.000000 2352.840000 2820.260000 2369.080000 ;
      RECT 0.000000 2352.420000 2819.520000 2352.840000 ;
      RECT 0.000000 2308.980000 2820.260000 2352.420000 ;
      RECT 0.740000 2308.560000 2820.260000 2308.980000 ;
      RECT 0.000000 2290.960000 2820.260000 2308.560000 ;
      RECT 0.000000 2290.540000 2819.520000 2290.960000 ;
      RECT 0.000000 2248.120000 2820.260000 2290.540000 ;
      RECT 0.740000 2247.700000 2820.260000 2248.120000 ;
      RECT 0.000000 2229.080000 2820.260000 2247.700000 ;
      RECT 0.000000 2228.660000 2819.520000 2229.080000 ;
      RECT 0.000000 2187.260000 2820.260000 2228.660000 ;
      RECT 0.740000 2186.840000 2820.260000 2187.260000 ;
      RECT 0.000000 2167.200000 2820.260000 2186.840000 ;
      RECT 0.000000 2166.780000 2819.520000 2167.200000 ;
      RECT 0.000000 2126.740000 2820.260000 2166.780000 ;
      RECT 0.740000 2126.320000 2820.260000 2126.740000 ;
      RECT 0.000000 2105.320000 2820.260000 2126.320000 ;
      RECT 0.000000 2104.900000 2819.520000 2105.320000 ;
      RECT 0.000000 2065.880000 2820.260000 2104.900000 ;
      RECT 0.740000 2065.460000 2820.260000 2065.880000 ;
      RECT 0.000000 2043.440000 2820.260000 2065.460000 ;
      RECT 0.000000 2043.020000 2819.520000 2043.440000 ;
      RECT 0.000000 2005.020000 2820.260000 2043.020000 ;
      RECT 0.740000 2004.600000 2820.260000 2005.020000 ;
      RECT 0.000000 1981.560000 2820.260000 2004.600000 ;
      RECT 0.000000 1981.140000 2819.520000 1981.560000 ;
      RECT 0.000000 1944.500000 2820.260000 1981.140000 ;
      RECT 0.740000 1944.080000 2820.260000 1944.500000 ;
      RECT 0.000000 1919.680000 2820.260000 1944.080000 ;
      RECT 0.000000 1919.260000 2819.520000 1919.680000 ;
      RECT 0.000000 1883.640000 2820.260000 1919.260000 ;
      RECT 0.740000 1883.220000 2820.260000 1883.640000 ;
      RECT 0.000000 1857.460000 2820.260000 1883.220000 ;
      RECT 0.000000 1857.040000 2819.520000 1857.460000 ;
      RECT 0.000000 1822.780000 2820.260000 1857.040000 ;
      RECT 0.740000 1822.360000 2820.260000 1822.780000 ;
      RECT 0.000000 1795.580000 2820.260000 1822.360000 ;
      RECT 0.000000 1795.160000 2819.520000 1795.580000 ;
      RECT 0.000000 1762.260000 2820.260000 1795.160000 ;
      RECT 0.740000 1761.840000 2820.260000 1762.260000 ;
      RECT 0.000000 1733.700000 2820.260000 1761.840000 ;
      RECT 0.000000 1733.280000 2819.520000 1733.700000 ;
      RECT 0.000000 1701.400000 2820.260000 1733.280000 ;
      RECT 0.740000 1700.980000 2820.260000 1701.400000 ;
      RECT 0.000000 1671.820000 2820.260000 1700.980000 ;
      RECT 0.000000 1671.400000 2819.520000 1671.820000 ;
      RECT 0.000000 1640.540000 2820.260000 1671.400000 ;
      RECT 0.740000 1640.120000 2820.260000 1640.540000 ;
      RECT 0.000000 1609.940000 2820.260000 1640.120000 ;
      RECT 0.000000 1609.520000 2819.520000 1609.940000 ;
      RECT 0.000000 1580.020000 2820.260000 1609.520000 ;
      RECT 0.740000 1579.600000 2820.260000 1580.020000 ;
      RECT 0.000000 1548.060000 2820.260000 1579.600000 ;
      RECT 0.000000 1547.640000 2819.520000 1548.060000 ;
      RECT 0.000000 1519.160000 2820.260000 1547.640000 ;
      RECT 0.740000 1518.740000 2820.260000 1519.160000 ;
      RECT 0.000000 1486.180000 2820.260000 1518.740000 ;
      RECT 0.000000 1485.760000 2819.520000 1486.180000 ;
      RECT 0.000000 1458.300000 2820.260000 1485.760000 ;
      RECT 0.740000 1457.880000 2820.260000 1458.300000 ;
      RECT 0.000000 1424.300000 2820.260000 1457.880000 ;
      RECT 0.000000 1423.880000 2819.520000 1424.300000 ;
      RECT 0.000000 1397.780000 2820.260000 1423.880000 ;
      RECT 0.740000 1397.360000 2820.260000 1397.780000 ;
      RECT 0.000000 1362.420000 2820.260000 1397.360000 ;
      RECT 0.000000 1362.000000 2819.520000 1362.420000 ;
      RECT 0.000000 1336.920000 2820.260000 1362.000000 ;
      RECT 0.740000 1336.500000 2820.260000 1336.920000 ;
      RECT 0.000000 1300.200000 2820.260000 1336.500000 ;
      RECT 0.000000 1299.780000 2819.520000 1300.200000 ;
      RECT 0.000000 1276.060000 2820.260000 1299.780000 ;
      RECT 0.740000 1275.640000 2820.260000 1276.060000 ;
      RECT 0.000000 1238.320000 2820.260000 1275.640000 ;
      RECT 0.000000 1237.900000 2819.520000 1238.320000 ;
      RECT 0.000000 1215.540000 2820.260000 1237.900000 ;
      RECT 0.740000 1215.120000 2820.260000 1215.540000 ;
      RECT 0.000000 1176.440000 2820.260000 1215.120000 ;
      RECT 0.000000 1176.020000 2819.520000 1176.440000 ;
      RECT 0.000000 1154.680000 2820.260000 1176.020000 ;
      RECT 0.740000 1154.260000 2820.260000 1154.680000 ;
      RECT 0.000000 1114.560000 2820.260000 1154.260000 ;
      RECT 0.000000 1114.140000 2819.520000 1114.560000 ;
      RECT 0.000000 1093.820000 2820.260000 1114.140000 ;
      RECT 0.740000 1093.400000 2820.260000 1093.820000 ;
      RECT 0.000000 1052.680000 2820.260000 1093.400000 ;
      RECT 0.000000 1052.260000 2819.520000 1052.680000 ;
      RECT 0.000000 1032.960000 2820.260000 1052.260000 ;
      RECT 0.740000 1032.540000 2820.260000 1032.960000 ;
      RECT 0.000000 990.800000 2820.260000 1032.540000 ;
      RECT 0.000000 990.380000 2819.520000 990.800000 ;
      RECT 0.000000 972.440000 2820.260000 990.380000 ;
      RECT 0.740000 972.020000 2820.260000 972.440000 ;
      RECT 0.000000 928.920000 2820.260000 972.020000 ;
      RECT 0.000000 928.500000 2819.520000 928.920000 ;
      RECT 0.000000 911.580000 2820.260000 928.500000 ;
      RECT 0.740000 911.160000 2820.260000 911.580000 ;
      RECT 0.000000 867.040000 2820.260000 911.160000 ;
      RECT 0.000000 866.620000 2819.520000 867.040000 ;
      RECT 0.000000 850.720000 2820.260000 866.620000 ;
      RECT 0.740000 850.300000 2820.260000 850.720000 ;
      RECT 0.000000 804.820000 2820.260000 850.300000 ;
      RECT 0.000000 804.400000 2819.520000 804.820000 ;
      RECT 0.000000 790.200000 2820.260000 804.400000 ;
      RECT 0.740000 789.780000 2820.260000 790.200000 ;
      RECT 0.000000 742.940000 2820.260000 789.780000 ;
      RECT 0.000000 742.520000 2819.520000 742.940000 ;
      RECT 0.000000 729.340000 2820.260000 742.520000 ;
      RECT 0.740000 728.920000 2820.260000 729.340000 ;
      RECT 0.000000 681.060000 2820.260000 728.920000 ;
      RECT 0.000000 680.640000 2819.520000 681.060000 ;
      RECT 0.000000 668.480000 2820.260000 680.640000 ;
      RECT 0.740000 668.060000 2820.260000 668.480000 ;
      RECT 0.000000 619.180000 2820.260000 668.060000 ;
      RECT 0.000000 618.760000 2819.520000 619.180000 ;
      RECT 0.000000 607.960000 2820.260000 618.760000 ;
      RECT 0.740000 607.540000 2820.260000 607.960000 ;
      RECT 0.000000 557.300000 2820.260000 607.540000 ;
      RECT 0.000000 556.880000 2819.520000 557.300000 ;
      RECT 0.000000 547.100000 2820.260000 556.880000 ;
      RECT 0.740000 546.680000 2820.260000 547.100000 ;
      RECT 0.000000 495.420000 2820.260000 546.680000 ;
      RECT 0.000000 495.000000 2819.520000 495.420000 ;
      RECT 0.000000 486.240000 2820.260000 495.000000 ;
      RECT 0.740000 485.820000 2820.260000 486.240000 ;
      RECT 0.000000 433.540000 2820.260000 485.820000 ;
      RECT 0.000000 433.120000 2819.520000 433.540000 ;
      RECT 0.000000 425.720000 2820.260000 433.120000 ;
      RECT 0.740000 425.300000 2820.260000 425.720000 ;
      RECT 0.000000 371.660000 2820.260000 425.300000 ;
      RECT 0.000000 371.240000 2819.520000 371.660000 ;
      RECT 0.000000 364.860000 2820.260000 371.240000 ;
      RECT 0.740000 364.440000 2820.260000 364.860000 ;
      RECT 0.000000 309.780000 2820.260000 364.440000 ;
      RECT 0.000000 309.360000 2819.520000 309.780000 ;
      RECT 0.000000 304.000000 2820.260000 309.360000 ;
      RECT 0.740000 303.580000 2820.260000 304.000000 ;
      RECT 0.000000 247.560000 2820.260000 303.580000 ;
      RECT 0.000000 247.140000 2819.520000 247.560000 ;
      RECT 0.000000 243.480000 2820.260000 247.140000 ;
      RECT 0.740000 243.060000 2820.260000 243.480000 ;
      RECT 0.000000 185.680000 2820.260000 243.060000 ;
      RECT 0.000000 185.260000 2819.520000 185.680000 ;
      RECT 0.000000 182.620000 2820.260000 185.260000 ;
      RECT 0.740000 182.200000 2820.260000 182.620000 ;
      RECT 0.000000 123.800000 2820.260000 182.200000 ;
      RECT 0.000000 123.380000 2819.520000 123.800000 ;
      RECT 0.000000 121.760000 2820.260000 123.380000 ;
      RECT 0.740000 121.340000 2820.260000 121.760000 ;
      RECT 0.000000 61.920000 2820.260000 121.340000 ;
      RECT 0.000000 61.500000 2819.520000 61.920000 ;
      RECT 0.000000 61.240000 2820.260000 61.500000 ;
      RECT 0.740000 60.820000 2820.260000 61.240000 ;
      RECT 0.000000 2.420000 2820.260000 60.820000 ;
      RECT 0.740000 2.080000 2820.260000 2.420000 ;
      RECT 0.740000 2.000000 2819.520000 2.080000 ;
      RECT 0.000000 1.660000 2819.520000 2.000000 ;
      RECT 0.000000 0.000000 2820.260000 1.660000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 2820.260000 3219.800000 ;
    LAYER met4 ;
      RECT 0.000000 1742.830000 2820.260000 3219.800000 ;
      RECT 4.460000 1732.130000 2820.260000 1742.830000 ;
      RECT 4.460000 1730.187000 5.660000 1732.130000 ;
      RECT 0.000000 1730.187000 1.860000 1742.830000 ;
      RECT 8.260000 1716.105000 2820.260000 1732.130000 ;
      RECT 0.000000 1716.105000 5.660000 1730.187000 ;
      RECT 0.000000 0.000000 2820.260000 1716.105000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2820.260000 3219.800000 ;
  END
END user_proj_example

END LIBRARY
