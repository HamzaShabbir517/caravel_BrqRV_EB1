module eb1_brqrv_wrapper (
`ifdef USE_POWER_PINS
	VPWR,
	VGND,
`endif	
	clk,
	rst_l,
	dbg_rst_l,
	rst_vec,
	nmi_int,
	nmi_vec,
	jtag_id,
	uart_rx,
	trace_rv_i_insn_ip,
	trace_rv_i_address_ip,
	trace_rv_i_valid_ip,
	trace_rv_i_exception_ip,
	trace_rv_i_ecause_ip,
	trace_rv_i_interrupt_ip,
	trace_rv_i_tval_ip,
	lsu_axi_awvalid,
	lsu_axi_awready,
	lsu_axi_awid,
	lsu_axi_awaddr,
	lsu_axi_awregion,
	lsu_axi_awlen,
	lsu_axi_awsize,
	lsu_axi_awburst,
	lsu_axi_awlock,
	lsu_axi_awcache,
	lsu_axi_awprot,
	lsu_axi_awqos,
	lsu_axi_wvalid,
	lsu_axi_wready,
	lsu_axi_wdata,
	lsu_axi_wstrb,
	lsu_axi_wlast,
	lsu_axi_bvalid,
	lsu_axi_bready,
	lsu_axi_bresp,
	lsu_axi_bid,
	lsu_axi_arvalid,
	lsu_axi_arready,
	lsu_axi_arid,
	lsu_axi_araddr,
	lsu_axi_arregion,
	lsu_axi_arlen,
	lsu_axi_arsize,
	lsu_axi_arburst,
	lsu_axi_arlock,
	lsu_axi_arcache,
	lsu_axi_arprot,
	lsu_axi_arqos,
	lsu_axi_rvalid,
	lsu_axi_rready,
	lsu_axi_rid,
	lsu_axi_rdata,
	lsu_axi_rresp,
	lsu_axi_rlast,
	ifu_axi_awvalid,
	ifu_axi_awready,
	ifu_axi_awid,
	ifu_axi_awaddr,
	ifu_axi_awregion,
	ifu_axi_awlen,
	ifu_axi_awsize,
	ifu_axi_awburst,
	ifu_axi_awlock,
	ifu_axi_awcache,
	ifu_axi_awprot,
	ifu_axi_awqos,
	ifu_axi_wvalid,
	ifu_axi_wready,
	ifu_axi_wdata,
	ifu_axi_wstrb,
	ifu_axi_wlast,
	ifu_axi_bvalid,
	ifu_axi_bready,
	ifu_axi_bresp,
	ifu_axi_bid,
	ifu_axi_arvalid,
	ifu_axi_arready,
	ifu_axi_arid,
	ifu_axi_araddr,
	ifu_axi_arregion,
	ifu_axi_arlen,
	ifu_axi_arsize,
	ifu_axi_arburst,
	ifu_axi_arlock,
	ifu_axi_arcache,
	ifu_axi_arprot,
	ifu_axi_arqos,
	ifu_axi_rvalid,
	ifu_axi_rready,
	ifu_axi_rid,
	ifu_axi_rdata,
	ifu_axi_rresp,
	ifu_axi_rlast,
	sb_axi_awvalid,
	sb_axi_awready,
	sb_axi_awid,
	sb_axi_awaddr,
	sb_axi_awregion,
	sb_axi_awlen,
	sb_axi_awsize,
	sb_axi_awburst,
	sb_axi_awlock,
	sb_axi_awcache,
	sb_axi_awprot,
	sb_axi_awqos,
	sb_axi_wvalid,
	sb_axi_wready,
	sb_axi_wdata,
	sb_axi_wstrb,
	sb_axi_wlast,
	sb_axi_bvalid,
	sb_axi_bready,
	sb_axi_bresp,
	sb_axi_bid,
	sb_axi_arvalid,
	sb_axi_arready,
	sb_axi_arid,
	sb_axi_araddr,
	sb_axi_arregion,
	sb_axi_arlen,
	sb_axi_arsize,
	sb_axi_arburst,
	sb_axi_arlock,
	sb_axi_arcache,
	sb_axi_arprot,
	sb_axi_arqos,
	sb_axi_rvalid,
	sb_axi_rready,
	sb_axi_rid,
	sb_axi_rdata,
	sb_axi_rresp,
	sb_axi_rlast,
	dma_axi_awvalid,
	dma_axi_awready,
	dma_axi_awid,
	dma_axi_awaddr,
	dma_axi_awsize,
	dma_axi_awprot,
	dma_axi_awlen,
	dma_axi_awburst,
	dma_axi_wvalid,
	dma_axi_wready,
	dma_axi_wdata,
	dma_axi_wstrb,
	dma_axi_wlast,
	dma_axi_bvalid,
	dma_axi_bready,
	dma_axi_bresp,
	dma_axi_bid,
	dma_axi_arvalid,
	dma_axi_arready,
	dma_axi_arid,
	dma_axi_araddr,
	dma_axi_arsize,
	dma_axi_arprot,
	dma_axi_arlen,
	dma_axi_arburst,
	dma_axi_rvalid,
	dma_axi_rready,
	dma_axi_rid,
	dma_axi_rdata,
	dma_axi_rresp,
	dma_axi_rlast,
	lsu_bus_clk_en,
	ifu_bus_clk_en,
	dbg_bus_clk_en,
	dma_bus_clk_en,
	dccm_ext_in_pkt,
	iccm_ext_in_pkt,
	ic_data_ext_in_pkt,
	ic_tag_ext_in_pkt,
	timer_int,
	soft_int,
	extintsrc_req,
	dec_tlu_perfcnt0,
	dec_tlu_perfcnt1,
	dec_tlu_perfcnt2,
	dec_tlu_perfcnt3,
	jtag_tck,
	jtag_tms,
	jtag_tdi,
	jtag_trst_n,
	jtag_tdo,
	core_id,
	mpc_debug_halt_req,
	mpc_debug_run_req,
	mpc_reset_run_req,
	mpc_debug_halt_ack,
	mpc_debug_run_ack,
	debug_brkpt_status,
	i_cpu_halt_req,
	o_cpu_halt_ack,
	o_cpu_halt_status,
	o_debug_mode_status,
	i_cpu_run_req,
	o_cpu_run_ack,
	scan_mode,
	mbist_mode,
	CLKS_PER_BIT
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
`ifdef USE_POWER_PINS
	inout wire VPWR;
	inout wire VGND;
`endif
	input wire clk;
	input wire rst_l;
	input wire dbg_rst_l;
	input wire [31:1] rst_vec;
	input wire nmi_int;
	input wire [31:1] nmi_vec;
	input wire [31:1] jtag_id;
	input uart_rx;
	output wire [31:0] trace_rv_i_insn_ip;
	output wire [31:0] trace_rv_i_address_ip;
	output wire trace_rv_i_valid_ip;
	output wire trace_rv_i_exception_ip;
	output wire [4:0] trace_rv_i_ecause_ip;
	output wire trace_rv_i_interrupt_ip;
	output wire [31:0] trace_rv_i_tval_ip;
	output wire lsu_axi_awvalid;
	input wire lsu_axi_awready;
	output wire [pt[181-:8] - 1:0] lsu_axi_awid;
	output wire [31:0] lsu_axi_awaddr;
	output wire [3:0] lsu_axi_awregion;
	output wire [7:0] lsu_axi_awlen;
	output wire [2:0] lsu_axi_awsize;
	output wire [1:0] lsu_axi_awburst;
	output wire lsu_axi_awlock;
	output wire [3:0] lsu_axi_awcache;
	output wire [2:0] lsu_axi_awprot;
	output wire [3:0] lsu_axi_awqos;
	output wire lsu_axi_wvalid;
	input wire lsu_axi_wready;
	output wire [63:0] lsu_axi_wdata;
	output wire [7:0] lsu_axi_wstrb;
	output wire lsu_axi_wlast;
	input wire lsu_axi_bvalid;
	output wire lsu_axi_bready;
	input wire [1:0] lsu_axi_bresp;
	input wire [pt[181-:8] - 1:0] lsu_axi_bid;
	output wire lsu_axi_arvalid;
	input wire lsu_axi_arready;
	output wire [pt[181-:8] - 1:0] lsu_axi_arid;
	output wire [31:0] lsu_axi_araddr;
	output wire [3:0] lsu_axi_arregion;
	output wire [7:0] lsu_axi_arlen;
	output wire [2:0] lsu_axi_arsize;
	output wire [1:0] lsu_axi_arburst;
	output wire lsu_axi_arlock;
	output wire [3:0] lsu_axi_arcache;
	output wire [2:0] lsu_axi_arprot;
	output wire [3:0] lsu_axi_arqos;
	input wire lsu_axi_rvalid;
	output wire lsu_axi_rready;
	input wire [pt[181-:8] - 1:0] lsu_axi_rid;
	input wire [63:0] lsu_axi_rdata;
	input wire [1:0] lsu_axi_rresp;
	input wire lsu_axi_rlast;
	output wire ifu_axi_awvalid;
	input wire ifu_axi_awready;
	output wire [pt[826-:8] - 1:0] ifu_axi_awid;
	output wire [31:0] ifu_axi_awaddr;
	output wire [3:0] ifu_axi_awregion;
	output wire [7:0] ifu_axi_awlen;
	output wire [2:0] ifu_axi_awsize;
	output wire [1:0] ifu_axi_awburst;
	output wire ifu_axi_awlock;
	output wire [3:0] ifu_axi_awcache;
	output wire [2:0] ifu_axi_awprot;
	output wire [3:0] ifu_axi_awqos;
	output wire ifu_axi_wvalid;
	input wire ifu_axi_wready;
	output wire [63:0] ifu_axi_wdata;
	output wire [7:0] ifu_axi_wstrb;
	output wire ifu_axi_wlast;
	input wire ifu_axi_bvalid;
	output wire ifu_axi_bready;
	input wire [1:0] ifu_axi_bresp;
	input wire [pt[826-:8] - 1:0] ifu_axi_bid;
	output wire ifu_axi_arvalid;
	input wire ifu_axi_arready;
	output wire [pt[826-:8] - 1:0] ifu_axi_arid;
	output wire [31:0] ifu_axi_araddr;
	output wire [3:0] ifu_axi_arregion;
	output wire [7:0] ifu_axi_arlen;
	output wire [2:0] ifu_axi_arsize;
	output wire [1:0] ifu_axi_arburst;
	output wire ifu_axi_arlock;
	output wire [3:0] ifu_axi_arcache;
	output wire [2:0] ifu_axi_arprot;
	output wire [3:0] ifu_axi_arqos;
	input wire ifu_axi_rvalid;
	output wire ifu_axi_rready;
	input wire [pt[826-:8] - 1:0] ifu_axi_rid;
	input wire [63:0] ifu_axi_rdata;
	input wire [1:0] ifu_axi_rresp;
	input wire ifu_axi_rlast;
	output wire sb_axi_awvalid;
	input wire sb_axi_awready;
	output wire [pt[12-:8] - 1:0] sb_axi_awid;
	output wire [31:0] sb_axi_awaddr;
	output wire [3:0] sb_axi_awregion;
	output wire [7:0] sb_axi_awlen;
	output wire [2:0] sb_axi_awsize;
	output wire [1:0] sb_axi_awburst;
	output wire sb_axi_awlock;
	output wire [3:0] sb_axi_awcache;
	output wire [2:0] sb_axi_awprot;
	output wire [3:0] sb_axi_awqos;
	output wire sb_axi_wvalid;
	input wire sb_axi_wready;
	output wire [63:0] sb_axi_wdata;
	output wire [7:0] sb_axi_wstrb;
	output wire sb_axi_wlast;
	input wire sb_axi_bvalid;
	output wire sb_axi_bready;
	input wire [1:0] sb_axi_bresp;
	input wire [pt[12-:8] - 1:0] sb_axi_bid;
	output wire sb_axi_arvalid;
	input wire sb_axi_arready;
	output wire [pt[12-:8] - 1:0] sb_axi_arid;
	output wire [31:0] sb_axi_araddr;
	output wire [3:0] sb_axi_arregion;
	output wire [7:0] sb_axi_arlen;
	output wire [2:0] sb_axi_arsize;
	output wire [1:0] sb_axi_arburst;
	output wire sb_axi_arlock;
	output wire [3:0] sb_axi_arcache;
	output wire [2:0] sb_axi_arprot;
	output wire [3:0] sb_axi_arqos;
	input wire sb_axi_rvalid;
	output wire sb_axi_rready;
	input wire [pt[12-:8] - 1:0] sb_axi_rid;
	input wire [63:0] sb_axi_rdata;
	input wire [1:0] sb_axi_rresp;
	input wire sb_axi_rlast;
	input wire dma_axi_awvalid;
	output wire dma_axi_awready;
	input wire [pt[1235-:8] - 1:0] dma_axi_awid;
	input wire [31:0] dma_axi_awaddr;
	input wire [2:0] dma_axi_awsize;
	input wire [2:0] dma_axi_awprot;
	input wire [7:0] dma_axi_awlen;
	input wire [1:0] dma_axi_awburst;
	input wire dma_axi_wvalid;
	output wire dma_axi_wready;
	input wire [63:0] dma_axi_wdata;
	input wire [7:0] dma_axi_wstrb;
	input wire dma_axi_wlast;
	output wire dma_axi_bvalid;
	input wire dma_axi_bready;
	output wire [1:0] dma_axi_bresp;
	output wire [pt[1235-:8] - 1:0] dma_axi_bid;
	input wire dma_axi_arvalid;
	output wire dma_axi_arready;
	input wire [pt[1235-:8] - 1:0] dma_axi_arid;
	input wire [31:0] dma_axi_araddr;
	input wire [2:0] dma_axi_arsize;
	input wire [2:0] dma_axi_arprot;
	input wire [7:0] dma_axi_arlen;
	input wire [1:0] dma_axi_arburst;
	output wire dma_axi_rvalid;
	input wire dma_axi_rready;
	output wire [pt[1235-:8] - 1:0] dma_axi_rid;
	output wire [63:0] dma_axi_rdata;
	output wire [1:0] dma_axi_rresp;
	output wire dma_axi_rlast;
	input wire lsu_bus_clk_en;
	input wire ifu_bus_clk_en;
	input wire dbg_bus_clk_en;
	input wire dma_bus_clk_en;
	input wire [(pt[1342-:9] * 12) - 1:0] dccm_ext_in_pkt;
	input wire [(pt[909-:9] * 12) - 1:0] iccm_ext_in_pkt;
	input wire [((pt[1060-:7] * pt[1189-:7]) * 12) - 1:0] ic_data_ext_in_pkt;
	input wire [(pt[1060-:7] * 12) - 1:0] ic_tag_ext_in_pkt;
	input wire timer_int;
	input wire soft_int;
	input wire [pt[56-:12]:1] extintsrc_req;
	output wire dec_tlu_perfcnt0;
	output wire dec_tlu_perfcnt1;
	output wire dec_tlu_perfcnt2;
	output wire dec_tlu_perfcnt3;
	input wire jtag_tck;
	input wire jtag_tms;
	input wire jtag_tdi;
	input wire jtag_trst_n;
	output wire jtag_tdo;
	input wire [31:4] core_id;
	input wire mpc_debug_halt_req;
	input wire mpc_debug_run_req;
	input wire mpc_reset_run_req;
	output wire mpc_debug_halt_ack;
	output wire mpc_debug_run_ack;
	output wire debug_brkpt_status;
	input wire i_cpu_halt_req;
	output wire o_cpu_halt_ack;
	output wire o_cpu_halt_status;
	output wire o_debug_mode_status;
	input wire i_cpu_run_req;
	output wire o_cpu_run_ack;
	input wire scan_mode;
	input wire mbist_mode;
	input [15:0] CLKS_PER_BIT;
	wire active_l2clk;
	wire free_l2clk;
	wire dccm_wren;
	wire dccm_rden;
	wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	wire [31:1] ic_rw_addr;
	wire [pt[1060-:7] - 1:0] ic_wr_en;
	wire ic_rd_en;
	wire [pt[1060-:7] - 1:0] ic_tag_valid;
	wire [pt[1060-:7] - 1:0] ic_rd_hit;
	wire ic_tag_perr;
	wire [pt[1104-:9]:3] ic_debug_addr;
	wire ic_debug_rd_en;
	wire ic_debug_wr_en;
	wire ic_debug_tag_array;
	wire [pt[1060-:7] - 1:0] ic_debug_way;
	wire [25:0] ictag_debug_rd_data;
	wire [(pt[1189-:7] * 71) - 1:0] ic_wr_data;
	wire [63:0] ic_rd_data;
	wire [70:0] ic_debug_rd_data;
	wire [70:0] ic_debug_wr_data;
	wire [pt[1189-:7] - 1:0] ic_eccerr;
	wire [pt[1189-:7] - 1:0] ic_parerr;
	wire [63:0] ic_premux_data;
	wire ic_sel_premux_data;
	wire [pt[936-:9] - 1:1] iccm_rw_addr;
	wire iccm_wren;
	wire iccm_rden;
	wire [2:0] iccm_wr_size;
	wire [77:0] iccm_wr_data;
	wire iccm_buf_correct_ecc;
	wire iccm_correction_state;
	wire [63:0] iccm_rd_data;
	wire [77:0] iccm_rd_data_ecc;
	wire core_rst;
	wire core_rst_l;
	wire jtag_tdoEn;
	wire dccm_clk_override;
	wire icm_clk_override;
	wire dec_tlu_core_ecc_disable;
	wire [31:0] haddr;
	wire [2:0] hburst;
	wire hmastlock;
	wire [3:0] hprot;
	wire [2:0] hsize;
	wire [1:0] htrans;
	wire hwrite;
	wire [63:0] hrdata;
	wire hready;
	wire hresp;
	wire [31:0] lsu_haddr;
	wire [2:0] lsu_hburst;
	wire lsu_hmastlock;
	wire [3:0] lsu_hprot;
	wire [2:0] lsu_hsize;
	wire [1:0] lsu_htrans;
	wire lsu_hwrite;
	wire [63:0] lsu_hwdata;
	wire [63:0] lsu_hrdata;
	wire lsu_hready;
	wire lsu_hresp;
	wire [31:0] sb_haddr;
	wire [2:0] sb_hburst;
	wire sb_hmastlock;
	wire [3:0] sb_hprot;
	wire [2:0] sb_hsize;
	wire [1:0] sb_htrans;
	wire sb_hwrite;
	wire [63:0] sb_hwdata;
	wire [63:0] sb_hrdata;
	wire sb_hready;
	wire sb_hresp;
	wire dma_hsel;
	wire [31:0] dma_haddr;
	wire [2:0] dma_hburst;
	wire dma_hmastlock;
	wire [3:0] dma_hprot;
	wire [2:0] dma_hsize;
	wire [1:0] dma_htrans;
	wire dma_hwrite;
	wire [63:0] dma_hwdata;
	wire dma_hreadyin;
	wire [63:0] dma_hrdata;
	wire dma_hreadyout;
	wire dma_hresp;
	assign hrdata[63:0] = {64 {1'sb0}};
	assign hready = 1'b0;
	assign hresp = 1'b0;
	assign lsu_hrdata[63:0] = {64 {1'sb0}};
	assign lsu_hready = 1'b0;
	assign lsu_hresp = 1'b0;
	assign sb_hrdata[63:0] = {64 {1'sb0}};
	assign sb_hready = 1'b0;
	assign sb_hresp = 1'b0;
	assign dma_hsel = 1'b0;
	assign dma_haddr[31:0] = {32 {1'sb0}};
	assign dma_hburst[2:0] = {3 {1'sb0}};
	assign dma_hmastlock = 1'b0;
	assign dma_hprot[3:0] = {4 {1'sb0}};
	assign dma_hsize[2:0] = {3 {1'sb0}};
	assign dma_htrans[1:0] = {2 {1'sb0}};
	assign dma_hwrite = 1'b0;
	assign dma_hwdata[63:0] = {64 {1'sb0}};
	assign dma_hreadyin = 1'b0;
	wire dmi_reg_en;
	wire [6:0] dmi_reg_addr;
	wire dmi_reg_wr_en;
	wire [31:0] dmi_reg_wdata;
	wire [31:0] dmi_reg_rdata;
	wire rx_dv_i;
	wire [7:0] rx_byte_i;
	wire iccm_instr_we;
	wire [13:0] iccm_instr_addr;
	wire [31:0] iccm_instr_wdata;
	eb1_brqrv #(.pt(pt)) brqrv(
		.clk(clk),
		.rst_l(core_rst),
		.dbg_rst_l(dbg_rst_l),
		.rst_vec(rst_vec),
		.nmi_int(nmi_int),
		.nmi_vec(nmi_vec),
		.core_rst_l(core_rst_l),
		.active_l2clk(active_l2clk),
		.free_l2clk(free_l2clk),
		.trace_rv_i_insn_ip(trace_rv_i_insn_ip),
		.trace_rv_i_address_ip(trace_rv_i_address_ip),
		.trace_rv_i_valid_ip(trace_rv_i_valid_ip),
		.trace_rv_i_exception_ip(trace_rv_i_exception_ip),
		.trace_rv_i_ecause_ip(trace_rv_i_ecause_ip),
		.trace_rv_i_interrupt_ip(trace_rv_i_interrupt_ip),
		.trace_rv_i_tval_ip(trace_rv_i_tval_ip),
		.dccm_clk_override(dccm_clk_override),
		.icm_clk_override(icm_clk_override),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.i_cpu_halt_req(i_cpu_halt_req),
		.i_cpu_run_req(i_cpu_run_req),
		.o_cpu_halt_ack(o_cpu_halt_ack),
		.o_cpu_halt_status(o_cpu_halt_status),
		.o_cpu_run_ack(o_cpu_run_ack),
		.o_debug_mode_status(o_debug_mode_status),
		.core_id(core_id),
		.mpc_debug_halt_req(mpc_debug_halt_req),
		.mpc_debug_run_req(mpc_debug_run_req),
		.mpc_reset_run_req(mpc_reset_run_req),
		.mpc_debug_halt_ack(mpc_debug_halt_ack),
		.mpc_debug_run_ack(mpc_debug_run_ack),
		.debug_brkpt_status(debug_brkpt_status),
		.dec_tlu_perfcnt0(dec_tlu_perfcnt0),
		.dec_tlu_perfcnt1(dec_tlu_perfcnt1),
		.dec_tlu_perfcnt2(dec_tlu_perfcnt2),
		.dec_tlu_perfcnt3(dec_tlu_perfcnt3),
		.dccm_wren(dccm_wren),
		.dccm_rden(dccm_rden),
		.dccm_wr_addr_lo(dccm_wr_addr_lo),
		.dccm_wr_addr_hi(dccm_wr_addr_hi),
		.dccm_rd_addr_lo(dccm_rd_addr_lo),
		.dccm_rd_addr_hi(dccm_rd_addr_hi),
		.dccm_wr_data_lo(dccm_wr_data_lo),
		.dccm_wr_data_hi(dccm_wr_data_hi),
		.dccm_rd_data_lo(dccm_rd_data_lo),
		.dccm_rd_data_hi(dccm_rd_data_hi),
		.iccm_rw_addr(iccm_rw_addr),
		.iccm_wren(iccm_wren),
		.iccm_rden(iccm_rden),
		.iccm_wr_size(iccm_wr_size),
		.iccm_wr_data(iccm_wr_data),
		.iccm_buf_correct_ecc(iccm_buf_correct_ecc),
		.iccm_correction_state(iccm_correction_state),
		.iccm_rd_data(iccm_rd_data),
		.iccm_rd_data_ecc(iccm_rd_data_ecc),
		.ic_rw_addr(ic_rw_addr),
		.ic_tag_valid(ic_tag_valid),
		.ic_wr_en(ic_wr_en),
		.ic_rd_en(ic_rd_en),
		.ic_wr_data(ic_wr_data),
		.ic_rd_data(ic_rd_data),
		.ic_debug_rd_data(ic_debug_rd_data),
		.ictag_debug_rd_data(ictag_debug_rd_data),
		.ic_debug_wr_data(ic_debug_wr_data),
		.ic_eccerr(ic_eccerr),
		.ic_parerr(ic_parerr),
		.ic_premux_data(ic_premux_data),
		.ic_sel_premux_data(ic_sel_premux_data),
		.ic_debug_addr(ic_debug_addr),
		.ic_debug_rd_en(ic_debug_rd_en),
		.ic_debug_wr_en(ic_debug_wr_en),
		.ic_debug_tag_array(ic_debug_tag_array),
		.ic_debug_way(ic_debug_way),
		.ic_rd_hit(ic_rd_hit),
		.ic_tag_perr(ic_tag_perr),
		.lsu_axi_awvalid(lsu_axi_awvalid),
		.lsu_axi_awready(lsu_axi_awready),
		.lsu_axi_awid(lsu_axi_awid),
		.lsu_axi_awaddr(lsu_axi_awaddr),
		.lsu_axi_awregion(lsu_axi_awregion),
		.lsu_axi_awlen(lsu_axi_awlen),
		.lsu_axi_awsize(lsu_axi_awsize),
		.lsu_axi_awburst(lsu_axi_awburst),
		.lsu_axi_awlock(lsu_axi_awlock),
		.lsu_axi_awcache(lsu_axi_awcache),
		.lsu_axi_awprot(lsu_axi_awprot),
		.lsu_axi_awqos(lsu_axi_awqos),
		.lsu_axi_wvalid(lsu_axi_wvalid),
		.lsu_axi_wready(lsu_axi_wready),
		.lsu_axi_wdata(lsu_axi_wdata),
		.lsu_axi_wstrb(lsu_axi_wstrb),
		.lsu_axi_wlast(lsu_axi_wlast),
		.lsu_axi_bvalid(lsu_axi_bvalid),
		.lsu_axi_bready(lsu_axi_bready),
		.lsu_axi_bresp(lsu_axi_bresp),
		.lsu_axi_bid(lsu_axi_bid),
		.lsu_axi_arvalid(lsu_axi_arvalid),
		.lsu_axi_arready(lsu_axi_arready),
		.lsu_axi_arid(lsu_axi_arid),
		.lsu_axi_araddr(lsu_axi_araddr),
		.lsu_axi_arregion(lsu_axi_arregion),
		.lsu_axi_arlen(lsu_axi_arlen),
		.lsu_axi_arsize(lsu_axi_arsize),
		.lsu_axi_arburst(lsu_axi_arburst),
		.lsu_axi_arlock(lsu_axi_arlock),
		.lsu_axi_arcache(lsu_axi_arcache),
		.lsu_axi_arprot(lsu_axi_arprot),
		.lsu_axi_arqos(lsu_axi_arqos),
		.lsu_axi_rvalid(lsu_axi_rvalid),
		.lsu_axi_rready(lsu_axi_rready),
		.lsu_axi_rid(lsu_axi_rid),
		.lsu_axi_rdata(lsu_axi_rdata),
		.lsu_axi_rresp(lsu_axi_rresp),
		.lsu_axi_rlast(lsu_axi_rlast),
		.ifu_axi_awvalid(ifu_axi_awvalid),
		.ifu_axi_awready(ifu_axi_awready),
		.ifu_axi_awid(ifu_axi_awid),
		.ifu_axi_awaddr(ifu_axi_awaddr),
		.ifu_axi_awregion(ifu_axi_awregion),
		.ifu_axi_awlen(ifu_axi_awlen),
		.ifu_axi_awsize(ifu_axi_awsize),
		.ifu_axi_awburst(ifu_axi_awburst),
		.ifu_axi_awlock(ifu_axi_awlock),
		.ifu_axi_awcache(ifu_axi_awcache),
		.ifu_axi_awprot(ifu_axi_awprot),
		.ifu_axi_awqos(ifu_axi_awqos),
		.ifu_axi_wvalid(ifu_axi_wvalid),
		.ifu_axi_wready(ifu_axi_wready),
		.ifu_axi_wdata(ifu_axi_wdata),
		.ifu_axi_wstrb(ifu_axi_wstrb),
		.ifu_axi_wlast(ifu_axi_wlast),
		.ifu_axi_bvalid(ifu_axi_bvalid),
		.ifu_axi_bready(ifu_axi_bready),
		.ifu_axi_bresp(ifu_axi_bresp),
		.ifu_axi_bid(ifu_axi_bid),
		.ifu_axi_arvalid(ifu_axi_arvalid),
		.ifu_axi_arready(ifu_axi_arready),
		.ifu_axi_arid(ifu_axi_arid),
		.ifu_axi_araddr(ifu_axi_araddr),
		.ifu_axi_arregion(ifu_axi_arregion),
		.ifu_axi_arlen(ifu_axi_arlen),
		.ifu_axi_arsize(ifu_axi_arsize),
		.ifu_axi_arburst(ifu_axi_arburst),
		.ifu_axi_arlock(ifu_axi_arlock),
		.ifu_axi_arcache(ifu_axi_arcache),
		.ifu_axi_arprot(ifu_axi_arprot),
		.ifu_axi_arqos(ifu_axi_arqos),
		.ifu_axi_rvalid(ifu_axi_rvalid),
		.ifu_axi_rready(ifu_axi_rready),
		.ifu_axi_rid(ifu_axi_rid),
		.ifu_axi_rdata(ifu_axi_rdata),
		.ifu_axi_rresp(ifu_axi_rresp),
		.ifu_axi_rlast(ifu_axi_rlast),
		.sb_axi_awvalid(sb_axi_awvalid),
		.sb_axi_awready(sb_axi_awready),
		.sb_axi_awid(sb_axi_awid),
		.sb_axi_awaddr(sb_axi_awaddr),
		.sb_axi_awregion(sb_axi_awregion),
		.sb_axi_awlen(sb_axi_awlen),
		.sb_axi_awsize(sb_axi_awsize),
		.sb_axi_awburst(sb_axi_awburst),
		.sb_axi_awlock(sb_axi_awlock),
		.sb_axi_awcache(sb_axi_awcache),
		.sb_axi_awprot(sb_axi_awprot),
		.sb_axi_awqos(sb_axi_awqos),
		.sb_axi_wvalid(sb_axi_wvalid),
		.sb_axi_wready(sb_axi_wready),
		.sb_axi_wdata(sb_axi_wdata),
		.sb_axi_wstrb(sb_axi_wstrb),
		.sb_axi_wlast(sb_axi_wlast),
		.sb_axi_bvalid(sb_axi_bvalid),
		.sb_axi_bready(sb_axi_bready),
		.sb_axi_bresp(sb_axi_bresp),
		.sb_axi_bid(sb_axi_bid),
		.sb_axi_arvalid(sb_axi_arvalid),
		.sb_axi_arready(sb_axi_arready),
		.sb_axi_arid(sb_axi_arid),
		.sb_axi_araddr(sb_axi_araddr),
		.sb_axi_arregion(sb_axi_arregion),
		.sb_axi_arlen(sb_axi_arlen),
		.sb_axi_arsize(sb_axi_arsize),
		.sb_axi_arburst(sb_axi_arburst),
		.sb_axi_arlock(sb_axi_arlock),
		.sb_axi_arcache(sb_axi_arcache),
		.sb_axi_arprot(sb_axi_arprot),
		.sb_axi_arqos(sb_axi_arqos),
		.sb_axi_rvalid(sb_axi_rvalid),
		.sb_axi_rready(sb_axi_rready),
		.sb_axi_rid(sb_axi_rid),
		.sb_axi_rdata(sb_axi_rdata),
		.sb_axi_rresp(sb_axi_rresp),
		.sb_axi_rlast(sb_axi_rlast),
		.dma_axi_awvalid(dma_axi_awvalid),
		.dma_axi_awready(dma_axi_awready),
		.dma_axi_awid(dma_axi_awid),
		.dma_axi_awaddr(dma_axi_awaddr),
		.dma_axi_awsize(dma_axi_awsize),
		.dma_axi_awprot(dma_axi_awprot),
		.dma_axi_awlen(dma_axi_awlen),
		.dma_axi_awburst(dma_axi_awburst),
		.dma_axi_wvalid(dma_axi_wvalid),
		.dma_axi_wready(dma_axi_wready),
		.dma_axi_wdata(dma_axi_wdata),
		.dma_axi_wstrb(dma_axi_wstrb),
		.dma_axi_wlast(dma_axi_wlast),
		.dma_axi_bvalid(dma_axi_bvalid),
		.dma_axi_bready(dma_axi_bready),
		.dma_axi_bresp(dma_axi_bresp),
		.dma_axi_bid(dma_axi_bid),
		.dma_axi_arvalid(dma_axi_arvalid),
		.dma_axi_arready(dma_axi_arready),
		.dma_axi_arid(dma_axi_arid),
		.dma_axi_araddr(dma_axi_araddr),
		.dma_axi_arsize(dma_axi_arsize),
		.dma_axi_arprot(dma_axi_arprot),
		.dma_axi_arlen(dma_axi_arlen),
		.dma_axi_arburst(dma_axi_arburst),
		.dma_axi_rvalid(dma_axi_rvalid),
		.dma_axi_rready(dma_axi_rready),
		.dma_axi_rid(dma_axi_rid),
		.dma_axi_rdata(dma_axi_rdata),
		.dma_axi_rresp(dma_axi_rresp),
		.dma_axi_rlast(dma_axi_rlast),
		.haddr(haddr),
		.hburst(hburst),
		.hmastlock(hmastlock),
		.hprot(hprot),
		.hsize(hsize),
		.htrans(htrans),
		.hwrite(hwrite),
		.hrdata(hrdata),
		.hready(hready),
		.hresp(hresp),
		.lsu_haddr(lsu_haddr),
		.lsu_hburst(lsu_hburst),
		.lsu_hmastlock(lsu_hmastlock),
		.lsu_hprot(lsu_hprot),
		.lsu_hsize(lsu_hsize),
		.lsu_htrans(lsu_htrans),
		.lsu_hwrite(lsu_hwrite),
		.lsu_hwdata(lsu_hwdata),
		.lsu_hrdata(lsu_hrdata),
		.lsu_hready(lsu_hready),
		.lsu_hresp(lsu_hresp),
		.sb_haddr(sb_haddr),
		.sb_hburst(sb_hburst),
		.sb_hmastlock(sb_hmastlock),
		.sb_hprot(sb_hprot),
		.sb_hsize(sb_hsize),
		.sb_htrans(sb_htrans),
		.sb_hwrite(sb_hwrite),
		.sb_hwdata(sb_hwdata),
		.sb_hrdata(sb_hrdata),
		.sb_hready(sb_hready),
		.sb_hresp(sb_hresp),
		.dma_hsel(dma_hsel),
		.dma_haddr(dma_haddr),
		.dma_hburst(dma_hburst),
		.dma_hmastlock(dma_hmastlock),
		.dma_hprot(dma_hprot),
		.dma_hsize(dma_hsize),
		.dma_htrans(dma_htrans),
		.dma_hwrite(dma_hwrite),
		.dma_hwdata(dma_hwdata),
		.dma_hreadyin(dma_hreadyin),
		.dma_hrdata(dma_hrdata),
		.dma_hreadyout(dma_hreadyout),
		.dma_hresp(dma_hresp),
		.lsu_bus_clk_en(lsu_bus_clk_en),
		.ifu_bus_clk_en(ifu_bus_clk_en),
		.dbg_bus_clk_en(dbg_bus_clk_en),
		.dma_bus_clk_en(dma_bus_clk_en),
		.dmi_reg_en(dmi_reg_en),
		.dmi_reg_addr(dmi_reg_addr),
		.dmi_reg_wr_en(dmi_reg_wr_en),
		.dmi_reg_wdata(dmi_reg_wdata),
		.dmi_reg_rdata(dmi_reg_rdata),
		.extintsrc_req(extintsrc_req),
		.timer_int(timer_int),
		.soft_int(soft_int),
		.scan_mode(scan_mode)
	);
	eb1_mem #(.pt(pt)) mem(
		.clk(active_l2clk),
		.rst_l(rst_l),
		.iccm_rw_addr((core_rst ? iccm_rw_addr : iccm_instr_addr[10:0])),
		.iccm_wren((core_rst ? iccm_wren : iccm_instr_we)),
		.iccm_wr_data((core_rst ? iccm_wr_data : {7'h00, iccm_instr_wdata, 7'h00, iccm_instr_wdata})),
		.iccm_wr_size((core_rst ? iccm_wr_size : 3'b010)),
		`ifdef USE_POWER_PINS
		.VPWR(VPWR),
		.VGND(VGND),
		`endif
		.dccm_clk_override(dccm_clk_override),
		.icm_clk_override(icm_clk_override),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.dccm_wren(dccm_wren),
		.dccm_rden(dccm_rden),
		.dccm_wr_addr_lo(dccm_wr_addr_lo),
		.dccm_wr_addr_hi(dccm_wr_addr_hi),
		.dccm_rd_addr_lo(dccm_rd_addr_lo),
		.dccm_rd_addr_hi(dccm_rd_addr_hi),
		.dccm_wr_data_lo(dccm_wr_data_lo),
		.dccm_wr_data_hi(dccm_wr_data_hi),
		.dccm_rd_data_lo(dccm_rd_data_lo),
		.dccm_rd_data_hi(dccm_rd_data_hi),
		.dccm_ext_in_pkt(dccm_ext_in_pkt),
		.iccm_ext_in_pkt(iccm_ext_in_pkt),
		.iccm_buf_correct_ecc(iccm_buf_correct_ecc),
		.iccm_correction_state(iccm_correction_state),
		.iccm_rden(iccm_rden),
		.iccm_rd_data(iccm_rd_data),
		.iccm_rd_data_ecc(iccm_rd_data_ecc),
		.ic_rw_addr(ic_rw_addr),
		.ic_tag_valid(ic_tag_valid),
		.ic_wr_en(ic_wr_en),
		.ic_rd_en(ic_rd_en),
		.ic_premux_data(ic_premux_data),
		.ic_sel_premux_data(ic_sel_premux_data),
		.ic_data_ext_in_pkt(ic_data_ext_in_pkt),
		.ic_tag_ext_in_pkt(ic_tag_ext_in_pkt),
		.ic_wr_data(ic_wr_data),
		.ic_debug_wr_data(ic_debug_wr_data),
		.ic_debug_rd_data(ic_debug_rd_data),
		.ic_debug_addr(ic_debug_addr),
		.ic_debug_rd_en(ic_debug_rd_en),
		.ic_debug_wr_en(ic_debug_wr_en),
		.ic_debug_tag_array(ic_debug_tag_array),
		.ic_debug_way(ic_debug_way),
		.ic_rd_data(ic_rd_data),
		.ictag_debug_rd_data(ictag_debug_rd_data),
		.ic_eccerr(ic_eccerr),
		.ic_parerr(ic_parerr),
		.ic_rd_hit(ic_rd_hit),
		.ic_tag_perr(ic_tag_perr),
		.scan_mode(scan_mode)
	);
	eb1_iccm_controller iccm_controller(
		.clk_i(clk),
		.rst_ni(rst_l),
		.rx_dv_i(rx_dv_i),
		.rx_byte_i(rx_byte_i),
		.we_o(iccm_instr_we),
		.addr_o(iccm_instr_addr),
		.wdata_o(iccm_instr_wdata),
		.reset_o(core_rst)
	);
	eb1_uart_rx_prog uart_rx_m(
		.i_Clock(clk),
		.rst_ni(rst_l),
		.i_Rx_Serial(uart_rx),
		.CLKS_PER_BIT(CLKS_PER_BIT),
		.o_Rx_DV(rx_dv_i),
		.o_Rx_Byte(rx_byte_i)
	);
	dmi_wrapper dmi_wrapper(
		.trst_n(jtag_trst_n),
		.tck(jtag_tck),
		.tms(jtag_tms),
		.tdi(jtag_tdi),
		.tdo(jtag_tdo),
		.tdoEnable(),
		.core_rst_n(dbg_rst_l),
		.core_clk(clk),
		.jtag_id(jtag_id),
		.rd_data(dmi_reg_rdata),
		.reg_wr_data(dmi_reg_wdata),
		.reg_wr_addr(dmi_reg_addr),
		.reg_en(dmi_reg_en),
		.reg_wr_en(dmi_reg_wr_en),
		.dmi_hard_reset()
	);
endmodule
module eb1_brqrv (
	clk,
	rst_l,
	dbg_rst_l,
	rst_vec,
	nmi_int,
	nmi_vec,
	core_rst_l,
	active_l2clk,
	free_l2clk,
	trace_rv_i_insn_ip,
	trace_rv_i_address_ip,
	trace_rv_i_valid_ip,
	trace_rv_i_exception_ip,
	trace_rv_i_ecause_ip,
	trace_rv_i_interrupt_ip,
	trace_rv_i_tval_ip,
	dccm_clk_override,
	icm_clk_override,
	dec_tlu_core_ecc_disable,
	i_cpu_halt_req,
	i_cpu_run_req,
	o_cpu_halt_ack,
	o_cpu_halt_status,
	o_cpu_run_ack,
	o_debug_mode_status,
	core_id,
	mpc_debug_halt_req,
	mpc_debug_run_req,
	mpc_reset_run_req,
	mpc_debug_halt_ack,
	mpc_debug_run_ack,
	debug_brkpt_status,
	dec_tlu_perfcnt0,
	dec_tlu_perfcnt1,
	dec_tlu_perfcnt2,
	dec_tlu_perfcnt3,
	dccm_wren,
	dccm_rden,
	dccm_wr_addr_lo,
	dccm_wr_addr_hi,
	dccm_rd_addr_lo,
	dccm_rd_addr_hi,
	dccm_wr_data_lo,
	dccm_wr_data_hi,
	dccm_rd_data_lo,
	dccm_rd_data_hi,
	iccm_rw_addr,
	iccm_wren,
	iccm_rden,
	iccm_wr_size,
	iccm_wr_data,
	iccm_buf_correct_ecc,
	iccm_correction_state,
	iccm_rd_data,
	iccm_rd_data_ecc,
	ic_rw_addr,
	ic_tag_valid,
	ic_wr_en,
	ic_rd_en,
	ic_wr_data,
	ic_rd_data,
	ic_debug_rd_data,
	ictag_debug_rd_data,
	ic_debug_wr_data,
	ic_eccerr,
	ic_parerr,
	ic_premux_data,
	ic_sel_premux_data,
	ic_debug_addr,
	ic_debug_rd_en,
	ic_debug_wr_en,
	ic_debug_tag_array,
	ic_debug_way,
	ic_rd_hit,
	ic_tag_perr,
	lsu_axi_awvalid,
	lsu_axi_awready,
	lsu_axi_awid,
	lsu_axi_awaddr,
	lsu_axi_awregion,
	lsu_axi_awlen,
	lsu_axi_awsize,
	lsu_axi_awburst,
	lsu_axi_awlock,
	lsu_axi_awcache,
	lsu_axi_awprot,
	lsu_axi_awqos,
	lsu_axi_wvalid,
	lsu_axi_wready,
	lsu_axi_wdata,
	lsu_axi_wstrb,
	lsu_axi_wlast,
	lsu_axi_bvalid,
	lsu_axi_bready,
	lsu_axi_bresp,
	lsu_axi_bid,
	lsu_axi_arvalid,
	lsu_axi_arready,
	lsu_axi_arid,
	lsu_axi_araddr,
	lsu_axi_arregion,
	lsu_axi_arlen,
	lsu_axi_arsize,
	lsu_axi_arburst,
	lsu_axi_arlock,
	lsu_axi_arcache,
	lsu_axi_arprot,
	lsu_axi_arqos,
	lsu_axi_rvalid,
	lsu_axi_rready,
	lsu_axi_rid,
	lsu_axi_rdata,
	lsu_axi_rresp,
	lsu_axi_rlast,
	ifu_axi_awvalid,
	ifu_axi_awready,
	ifu_axi_awid,
	ifu_axi_awaddr,
	ifu_axi_awregion,
	ifu_axi_awlen,
	ifu_axi_awsize,
	ifu_axi_awburst,
	ifu_axi_awlock,
	ifu_axi_awcache,
	ifu_axi_awprot,
	ifu_axi_awqos,
	ifu_axi_wvalid,
	ifu_axi_wready,
	ifu_axi_wdata,
	ifu_axi_wstrb,
	ifu_axi_wlast,
	ifu_axi_bvalid,
	ifu_axi_bready,
	ifu_axi_bresp,
	ifu_axi_bid,
	ifu_axi_arvalid,
	ifu_axi_arready,
	ifu_axi_arid,
	ifu_axi_araddr,
	ifu_axi_arregion,
	ifu_axi_arlen,
	ifu_axi_arsize,
	ifu_axi_arburst,
	ifu_axi_arlock,
	ifu_axi_arcache,
	ifu_axi_arprot,
	ifu_axi_arqos,
	ifu_axi_rvalid,
	ifu_axi_rready,
	ifu_axi_rid,
	ifu_axi_rdata,
	ifu_axi_rresp,
	ifu_axi_rlast,
	sb_axi_awvalid,
	sb_axi_awready,
	sb_axi_awid,
	sb_axi_awaddr,
	sb_axi_awregion,
	sb_axi_awlen,
	sb_axi_awsize,
	sb_axi_awburst,
	sb_axi_awlock,
	sb_axi_awcache,
	sb_axi_awprot,
	sb_axi_awqos,
	sb_axi_wvalid,
	sb_axi_wready,
	sb_axi_wdata,
	sb_axi_wstrb,
	sb_axi_wlast,
	sb_axi_bvalid,
	sb_axi_bready,
	sb_axi_bresp,
	sb_axi_bid,
	sb_axi_arvalid,
	sb_axi_arready,
	sb_axi_arid,
	sb_axi_araddr,
	sb_axi_arregion,
	sb_axi_arlen,
	sb_axi_arsize,
	sb_axi_arburst,
	sb_axi_arlock,
	sb_axi_arcache,
	sb_axi_arprot,
	sb_axi_arqos,
	sb_axi_rvalid,
	sb_axi_rready,
	sb_axi_rid,
	sb_axi_rdata,
	sb_axi_rresp,
	sb_axi_rlast,
	dma_axi_awvalid,
	dma_axi_awready,
	dma_axi_awid,
	dma_axi_awaddr,
	dma_axi_awsize,
	dma_axi_awprot,
	dma_axi_awlen,
	dma_axi_awburst,
	dma_axi_wvalid,
	dma_axi_wready,
	dma_axi_wdata,
	dma_axi_wstrb,
	dma_axi_wlast,
	dma_axi_bvalid,
	dma_axi_bready,
	dma_axi_bresp,
	dma_axi_bid,
	dma_axi_arvalid,
	dma_axi_arready,
	dma_axi_arid,
	dma_axi_araddr,
	dma_axi_arsize,
	dma_axi_arprot,
	dma_axi_arlen,
	dma_axi_arburst,
	dma_axi_rvalid,
	dma_axi_rready,
	dma_axi_rid,
	dma_axi_rdata,
	dma_axi_rresp,
	dma_axi_rlast,
	haddr,
	hburst,
	hmastlock,
	hprot,
	hsize,
	htrans,
	hwrite,
	hrdata,
	hready,
	hresp,
	lsu_haddr,
	lsu_hburst,
	lsu_hmastlock,
	lsu_hprot,
	lsu_hsize,
	lsu_htrans,
	lsu_hwrite,
	lsu_hwdata,
	lsu_hrdata,
	lsu_hready,
	lsu_hresp,
	sb_haddr,
	sb_hburst,
	sb_hmastlock,
	sb_hprot,
	sb_hsize,
	sb_htrans,
	sb_hwrite,
	sb_hwdata,
	sb_hrdata,
	sb_hready,
	sb_hresp,
	dma_hsel,
	dma_haddr,
	dma_hburst,
	dma_hmastlock,
	dma_hprot,
	dma_hsize,
	dma_htrans,
	dma_hwrite,
	dma_hwdata,
	dma_hreadyin,
	dma_hrdata,
	dma_hreadyout,
	dma_hresp,
	lsu_bus_clk_en,
	ifu_bus_clk_en,
	dbg_bus_clk_en,
	dma_bus_clk_en,
	dmi_reg_en,
	dmi_reg_addr,
	dmi_reg_wr_en,
	dmi_reg_wdata,
	dmi_reg_rdata,
	extintsrc_req,
	timer_int,
	soft_int,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire dbg_rst_l;
	input wire [31:1] rst_vec;
	input wire nmi_int;
	input wire [31:1] nmi_vec;
	output wire core_rst_l;
	output wire active_l2clk;
	output wire free_l2clk;
	output wire [31:0] trace_rv_i_insn_ip;
	output wire [31:0] trace_rv_i_address_ip;
	output wire trace_rv_i_valid_ip;
	output wire trace_rv_i_exception_ip;
	output wire [4:0] trace_rv_i_ecause_ip;
	output wire trace_rv_i_interrupt_ip;
	output wire [31:0] trace_rv_i_tval_ip;
	output wire dccm_clk_override;
	output wire icm_clk_override;
	output wire dec_tlu_core_ecc_disable;
	input wire i_cpu_halt_req;
	input wire i_cpu_run_req;
	output wire o_cpu_halt_ack;
	output wire o_cpu_halt_status;
	output wire o_cpu_run_ack;
	output wire o_debug_mode_status;
	input wire [31:4] core_id;
	input wire mpc_debug_halt_req;
	input wire mpc_debug_run_req;
	input wire mpc_reset_run_req;
	output wire mpc_debug_halt_ack;
	output wire mpc_debug_run_ack;
	output wire debug_brkpt_status;
	output wire dec_tlu_perfcnt0;
	output wire dec_tlu_perfcnt1;
	output wire dec_tlu_perfcnt2;
	output wire dec_tlu_perfcnt3;
	output wire dccm_wren;
	output wire dccm_rden;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	output wire [pt[936-:9] - 1:1] iccm_rw_addr;
	output wire iccm_wren;
	output wire iccm_rden;
	output wire [2:0] iccm_wr_size;
	output wire [77:0] iccm_wr_data;
	output wire iccm_buf_correct_ecc;
	output wire iccm_correction_state;
	input wire [63:0] iccm_rd_data;
	input wire [77:0] iccm_rd_data_ecc;
	output wire [31:1] ic_rw_addr;
	output wire [pt[1060-:7] - 1:0] ic_tag_valid;
	output wire [pt[1060-:7] - 1:0] ic_wr_en;
	output wire ic_rd_en;
	output wire [(pt[1189-:7] * 71) - 1:0] ic_wr_data;
	input wire [63:0] ic_rd_data;
	input wire [70:0] ic_debug_rd_data;
	input wire [25:0] ictag_debug_rd_data;
	output wire [70:0] ic_debug_wr_data;
	input wire [pt[1189-:7] - 1:0] ic_eccerr;
	input wire [pt[1189-:7] - 1:0] ic_parerr;
	output wire [63:0] ic_premux_data;
	output wire ic_sel_premux_data;
	output wire [pt[1104-:9]:3] ic_debug_addr;
	output wire ic_debug_rd_en;
	output wire ic_debug_wr_en;
	output wire ic_debug_tag_array;
	output wire [pt[1060-:7] - 1:0] ic_debug_way;
	input wire [pt[1060-:7] - 1:0] ic_rd_hit;
	input wire ic_tag_perr;
	output wire lsu_axi_awvalid;
	input wire lsu_axi_awready;
	output wire [pt[181-:8] - 1:0] lsu_axi_awid;
	output wire [31:0] lsu_axi_awaddr;
	output wire [3:0] lsu_axi_awregion;
	output wire [7:0] lsu_axi_awlen;
	output wire [2:0] lsu_axi_awsize;
	output wire [1:0] lsu_axi_awburst;
	output wire lsu_axi_awlock;
	output wire [3:0] lsu_axi_awcache;
	output wire [2:0] lsu_axi_awprot;
	output wire [3:0] lsu_axi_awqos;
	output wire lsu_axi_wvalid;
	input wire lsu_axi_wready;
	output wire [63:0] lsu_axi_wdata;
	output wire [7:0] lsu_axi_wstrb;
	output wire lsu_axi_wlast;
	input wire lsu_axi_bvalid;
	output wire lsu_axi_bready;
	input wire [1:0] lsu_axi_bresp;
	input wire [pt[181-:8] - 1:0] lsu_axi_bid;
	output wire lsu_axi_arvalid;
	input wire lsu_axi_arready;
	output wire [pt[181-:8] - 1:0] lsu_axi_arid;
	output wire [31:0] lsu_axi_araddr;
	output wire [3:0] lsu_axi_arregion;
	output wire [7:0] lsu_axi_arlen;
	output wire [2:0] lsu_axi_arsize;
	output wire [1:0] lsu_axi_arburst;
	output wire lsu_axi_arlock;
	output wire [3:0] lsu_axi_arcache;
	output wire [2:0] lsu_axi_arprot;
	output wire [3:0] lsu_axi_arqos;
	input wire lsu_axi_rvalid;
	output wire lsu_axi_rready;
	input wire [pt[181-:8] - 1:0] lsu_axi_rid;
	input wire [63:0] lsu_axi_rdata;
	input wire [1:0] lsu_axi_rresp;
	input wire lsu_axi_rlast;
	output wire ifu_axi_awvalid;
	input wire ifu_axi_awready;
	output wire [pt[826-:8] - 1:0] ifu_axi_awid;
	output wire [31:0] ifu_axi_awaddr;
	output wire [3:0] ifu_axi_awregion;
	output wire [7:0] ifu_axi_awlen;
	output wire [2:0] ifu_axi_awsize;
	output wire [1:0] ifu_axi_awburst;
	output wire ifu_axi_awlock;
	output wire [3:0] ifu_axi_awcache;
	output wire [2:0] ifu_axi_awprot;
	output wire [3:0] ifu_axi_awqos;
	output wire ifu_axi_wvalid;
	input wire ifu_axi_wready;
	output wire [63:0] ifu_axi_wdata;
	output wire [7:0] ifu_axi_wstrb;
	output wire ifu_axi_wlast;
	input wire ifu_axi_bvalid;
	output wire ifu_axi_bready;
	input wire [1:0] ifu_axi_bresp;
	input wire [pt[826-:8] - 1:0] ifu_axi_bid;
	output wire ifu_axi_arvalid;
	input wire ifu_axi_arready;
	output wire [pt[826-:8] - 1:0] ifu_axi_arid;
	output wire [31:0] ifu_axi_araddr;
	output wire [3:0] ifu_axi_arregion;
	output wire [7:0] ifu_axi_arlen;
	output wire [2:0] ifu_axi_arsize;
	output wire [1:0] ifu_axi_arburst;
	output wire ifu_axi_arlock;
	output wire [3:0] ifu_axi_arcache;
	output wire [2:0] ifu_axi_arprot;
	output wire [3:0] ifu_axi_arqos;
	input wire ifu_axi_rvalid;
	output wire ifu_axi_rready;
	input wire [pt[826-:8] - 1:0] ifu_axi_rid;
	input wire [63:0] ifu_axi_rdata;
	input wire [1:0] ifu_axi_rresp;
	input wire ifu_axi_rlast;
	output wire sb_axi_awvalid;
	input wire sb_axi_awready;
	output wire [pt[12-:8] - 1:0] sb_axi_awid;
	output wire [31:0] sb_axi_awaddr;
	output wire [3:0] sb_axi_awregion;
	output wire [7:0] sb_axi_awlen;
	output wire [2:0] sb_axi_awsize;
	output wire [1:0] sb_axi_awburst;
	output wire sb_axi_awlock;
	output wire [3:0] sb_axi_awcache;
	output wire [2:0] sb_axi_awprot;
	output wire [3:0] sb_axi_awqos;
	output wire sb_axi_wvalid;
	input wire sb_axi_wready;
	output wire [63:0] sb_axi_wdata;
	output wire [7:0] sb_axi_wstrb;
	output wire sb_axi_wlast;
	input wire sb_axi_bvalid;
	output wire sb_axi_bready;
	input wire [1:0] sb_axi_bresp;
	input wire [pt[12-:8] - 1:0] sb_axi_bid;
	output wire sb_axi_arvalid;
	input wire sb_axi_arready;
	output wire [pt[12-:8] - 1:0] sb_axi_arid;
	output wire [31:0] sb_axi_araddr;
	output wire [3:0] sb_axi_arregion;
	output wire [7:0] sb_axi_arlen;
	output wire [2:0] sb_axi_arsize;
	output wire [1:0] sb_axi_arburst;
	output wire sb_axi_arlock;
	output wire [3:0] sb_axi_arcache;
	output wire [2:0] sb_axi_arprot;
	output wire [3:0] sb_axi_arqos;
	input wire sb_axi_rvalid;
	output wire sb_axi_rready;
	input wire [pt[12-:8] - 1:0] sb_axi_rid;
	input wire [63:0] sb_axi_rdata;
	input wire [1:0] sb_axi_rresp;
	input wire sb_axi_rlast;
	input wire dma_axi_awvalid;
	output wire dma_axi_awready;
	input wire [pt[1235-:8] - 1:0] dma_axi_awid;
	input wire [31:0] dma_axi_awaddr;
	input wire [2:0] dma_axi_awsize;
	input wire [2:0] dma_axi_awprot;
	input wire [7:0] dma_axi_awlen;
	input wire [1:0] dma_axi_awburst;
	input wire dma_axi_wvalid;
	output wire dma_axi_wready;
	input wire [63:0] dma_axi_wdata;
	input wire [7:0] dma_axi_wstrb;
	input wire dma_axi_wlast;
	output wire dma_axi_bvalid;
	input wire dma_axi_bready;
	output wire [1:0] dma_axi_bresp;
	output wire [pt[1235-:8] - 1:0] dma_axi_bid;
	input wire dma_axi_arvalid;
	output wire dma_axi_arready;
	input wire [pt[1235-:8] - 1:0] dma_axi_arid;
	input wire [31:0] dma_axi_araddr;
	input wire [2:0] dma_axi_arsize;
	input wire [2:0] dma_axi_arprot;
	input wire [7:0] dma_axi_arlen;
	input wire [1:0] dma_axi_arburst;
	output wire dma_axi_rvalid;
	input wire dma_axi_rready;
	output wire [pt[1235-:8] - 1:0] dma_axi_rid;
	output wire [63:0] dma_axi_rdata;
	output wire [1:0] dma_axi_rresp;
	output wire dma_axi_rlast;
	output wire [31:0] haddr;
	output wire [2:0] hburst;
	output wire hmastlock;
	output wire [3:0] hprot;
	output wire [2:0] hsize;
	output wire [1:0] htrans;
	output wire hwrite;
	input wire [63:0] hrdata;
	input wire hready;
	input wire hresp;
	output wire [31:0] lsu_haddr;
	output wire [2:0] lsu_hburst;
	output wire lsu_hmastlock;
	output wire [3:0] lsu_hprot;
	output wire [2:0] lsu_hsize;
	output wire [1:0] lsu_htrans;
	output wire lsu_hwrite;
	output wire [63:0] lsu_hwdata;
	input wire [63:0] lsu_hrdata;
	input wire lsu_hready;
	input wire lsu_hresp;
	output wire [31:0] sb_haddr;
	output wire [2:0] sb_hburst;
	output wire sb_hmastlock;
	output wire [3:0] sb_hprot;
	output wire [2:0] sb_hsize;
	output wire [1:0] sb_htrans;
	output wire sb_hwrite;
	output wire [63:0] sb_hwdata;
	input wire [63:0] sb_hrdata;
	input wire sb_hready;
	input wire sb_hresp;
	input wire dma_hsel;
	input wire [31:0] dma_haddr;
	input wire [2:0] dma_hburst;
	input wire dma_hmastlock;
	input wire [3:0] dma_hprot;
	input wire [2:0] dma_hsize;
	input wire [1:0] dma_htrans;
	input wire dma_hwrite;
	input wire [63:0] dma_hwdata;
	input wire dma_hreadyin;
	output wire [63:0] dma_hrdata;
	output wire dma_hreadyout;
	output wire dma_hresp;
	input wire lsu_bus_clk_en;
	input wire ifu_bus_clk_en;
	input wire dbg_bus_clk_en;
	input wire dma_bus_clk_en;
	input wire dmi_reg_en;
	input wire [6:0] dmi_reg_addr;
	input wire dmi_reg_wr_en;
	input wire [31:0] dmi_reg_wdata;
	output wire [31:0] dmi_reg_rdata;
	input wire [pt[56-:12]:1] extintsrc_req;
	input wire timer_int;
	input wire soft_int;
	input wire scan_mode;
	wire [63:0] hwdata_nc;
	wire ifu_pmu_instr_aligned;
	wire ifu_ic_error_start;
	wire ifu_iccm_rd_ecc_single_err;
	wire lsu_axi_awready_ahb;
	wire lsu_axi_wready_ahb;
	wire lsu_axi_bvalid_ahb;
	wire lsu_axi_bready_ahb;
	wire [1:0] lsu_axi_bresp_ahb;
	wire [pt[181-:8] - 1:0] lsu_axi_bid_ahb;
	wire lsu_axi_arready_ahb;
	wire lsu_axi_rvalid_ahb;
	wire [pt[181-:8] - 1:0] lsu_axi_rid_ahb;
	wire [63:0] lsu_axi_rdata_ahb;
	wire [1:0] lsu_axi_rresp_ahb;
	wire lsu_axi_rlast_ahb;
	wire lsu_axi_awready_int;
	wire lsu_axi_wready_int;
	wire lsu_axi_bvalid_int;
	wire lsu_axi_bready_int;
	wire [1:0] lsu_axi_bresp_int;
	wire [pt[181-:8] - 1:0] lsu_axi_bid_int;
	wire lsu_axi_arready_int;
	wire lsu_axi_rvalid_int;
	wire [pt[181-:8] - 1:0] lsu_axi_rid_int;
	wire [63:0] lsu_axi_rdata_int;
	wire [1:0] lsu_axi_rresp_int;
	wire lsu_axi_rlast_int;
	wire ifu_axi_awready_ahb;
	wire ifu_axi_wready_ahb;
	wire ifu_axi_bvalid_ahb;
	wire ifu_axi_bready_ahb;
	wire [1:0] ifu_axi_bresp_ahb;
	wire [pt[826-:8] - 1:0] ifu_axi_bid_ahb;
	wire ifu_axi_arready_ahb;
	wire ifu_axi_rvalid_ahb;
	wire [pt[826-:8] - 1:0] ifu_axi_rid_ahb;
	wire [63:0] ifu_axi_rdata_ahb;
	wire [1:0] ifu_axi_rresp_ahb;
	wire ifu_axi_rlast_ahb;
	wire ifu_axi_awready_int;
	wire ifu_axi_wready_int;
	wire ifu_axi_bvalid_int;
	wire ifu_axi_bready_int;
	wire [1:0] ifu_axi_bresp_int;
	wire [pt[826-:8] - 1:0] ifu_axi_bid_int;
	wire ifu_axi_arready_int;
	wire ifu_axi_rvalid_int;
	wire [pt[826-:8] - 1:0] ifu_axi_rid_int;
	wire [63:0] ifu_axi_rdata_int;
	wire [1:0] ifu_axi_rresp_int;
	wire ifu_axi_rlast_int;
	wire sb_axi_awready_ahb;
	wire sb_axi_wready_ahb;
	wire sb_axi_bvalid_ahb;
	wire sb_axi_bready_ahb;
	wire [1:0] sb_axi_bresp_ahb;
	wire [pt[12-:8] - 1:0] sb_axi_bid_ahb;
	wire sb_axi_arready_ahb;
	wire sb_axi_rvalid_ahb;
	wire [pt[12-:8] - 1:0] sb_axi_rid_ahb;
	wire [63:0] sb_axi_rdata_ahb;
	wire [1:0] sb_axi_rresp_ahb;
	wire sb_axi_rlast_ahb;
	wire sb_axi_awready_int;
	wire sb_axi_wready_int;
	wire sb_axi_bvalid_int;
	wire sb_axi_bready_int;
	wire [1:0] sb_axi_bresp_int;
	wire [pt[12-:8] - 1:0] sb_axi_bid_int;
	wire sb_axi_arready_int;
	wire sb_axi_rvalid_int;
	wire [pt[12-:8] - 1:0] sb_axi_rid_int;
	wire [63:0] sb_axi_rdata_int;
	wire [1:0] sb_axi_rresp_int;
	wire sb_axi_rlast_int;
	wire dma_axi_awvalid_ahb;
	wire [pt[1235-:8] - 1:0] dma_axi_awid_ahb;
	wire [31:0] dma_axi_awaddr_ahb;
	wire [2:0] dma_axi_awsize_ahb;
	wire [2:0] dma_axi_awprot_ahb;
	wire [7:0] dma_axi_awlen_ahb;
	wire [1:0] dma_axi_awburst_ahb;
	wire dma_axi_wvalid_ahb;
	wire [63:0] dma_axi_wdata_ahb;
	wire [7:0] dma_axi_wstrb_ahb;
	wire dma_axi_wlast_ahb;
	wire dma_axi_bready_ahb;
	wire dma_axi_arvalid_ahb;
	wire [pt[1235-:8] - 1:0] dma_axi_arid_ahb;
	wire [31:0] dma_axi_araddr_ahb;
	wire [2:0] dma_axi_arsize_ahb;
	wire [2:0] dma_axi_arprot_ahb;
	wire [7:0] dma_axi_arlen_ahb;
	wire [1:0] dma_axi_arburst_ahb;
	wire dma_axi_rready_ahb;
	wire dma_axi_awvalid_int;
	wire [pt[1235-:8] - 1:0] dma_axi_awid_int;
	wire [31:0] dma_axi_awaddr_int;
	wire [2:0] dma_axi_awsize_int;
	wire [2:0] dma_axi_awprot_int;
	wire [7:0] dma_axi_awlen_int;
	wire [1:0] dma_axi_awburst_int;
	wire dma_axi_wvalid_int;
	wire [63:0] dma_axi_wdata_int;
	wire [7:0] dma_axi_wstrb_int;
	wire dma_axi_wlast_int;
	wire dma_axi_bready_int;
	wire dma_axi_arvalid_int;
	wire [pt[1235-:8] - 1:0] dma_axi_arid_int;
	wire [31:0] dma_axi_araddr_int;
	wire [2:0] dma_axi_arsize_int;
	wire [2:0] dma_axi_arprot_int;
	wire [7:0] dma_axi_arlen_int;
	wire [1:0] dma_axi_arburst_int;
	wire dma_axi_rready_int;
	wire [70:0] ifu_ic_debug_rd_data;
	wire ifu_ic_debug_rd_data_valid;
	wire [89:0] dec_tlu_ic_diag_pkt;
	wire dec_i0_rs1_en_d;
	wire dec_i0_rs2_en_d;
	wire [31:0] gpr_i0_rs1_d;
	wire [31:0] gpr_i0_rs2_d;
	wire [31:0] dec_i0_result_r;
	wire [31:0] exu_i0_result_x;
	wire [31:1] exu_i0_pc_x;
	wire [31:1] exu_npc_r;
	wire [43:0] i0_ap;
	wire [151:0] trigger_pkt_any;
	wire [3:0] lsu_trigger_match_m;
	wire [31:0] dec_i0_immed_d;
	wire [12:1] dec_i0_br_immed_d;
	wire dec_i0_select_pc_d;
	wire [31:1] dec_i0_pc_d;
	wire [3:0] dec_i0_rs1_bypass_en_d;
	wire [3:0] dec_i0_rs2_bypass_en_d;
	wire dec_i0_alu_decode_d;
	wire dec_i0_branch_d;
	wire ifu_miss_state_idle;
	wire dec_tlu_flush_noredir_r;
	wire dec_tlu_flush_leak_one_r;
	wire dec_tlu_flush_err_r;
	wire ifu_i0_valid;
	wire [31:0] ifu_i0_instr;
	wire [31:1] ifu_i0_pc;
	wire exu_flush_final;
	wire [31:1] exu_flush_path_final;
	wire [31:0] exu_lsu_rs1_d;
	wire [31:0] exu_lsu_rs2_d;
	wire [13:0] lsu_p;
	wire dec_qual_lsu_d;
	wire dec_lsu_valid_raw_d;
	wire [11:0] dec_lsu_offset_d;
	wire [31:0] lsu_result_m;
	wire [31:0] lsu_result_corr_r;
	wire lsu_single_ecc_error_incr;
	wire [39:0] lsu_error_pkt_r;
	wire lsu_imprecise_error_load_any;
	wire lsu_imprecise_error_store_any;
	wire [31:0] lsu_imprecise_error_addr_any;
	wire lsu_load_stall_any;
	wire lsu_store_stall_any;
	wire lsu_idle_any;
	wire lsu_active;
	wire [31:1] lsu_fir_addr;
	wire [1:0] lsu_fir_error;
	wire lsu_nonblock_load_valid_m;
	wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	wire lsu_nonblock_load_inv_r;
	wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	wire lsu_nonblock_load_data_valid;
	wire [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	wire [31:0] lsu_nonblock_load_data;
	wire dec_csr_ren_d;
	wire [31:0] dec_csr_rddata_d;
	wire [31:0] exu_csr_rs1_x;
	wire dec_tlu_i0_commit_cmt;
	wire dec_tlu_flush_lower_r;
	wire dec_tlu_flush_lower_wb;
	wire dec_tlu_i0_kill_writeb_r;
	wire dec_tlu_fence_i_r;
	wire [31:1] dec_tlu_flush_path_r;
	wire [31:0] dec_tlu_mrac_ff;
	wire ifu_i0_pc4;
	wire [19:0] mul_p;
	wire [2:0] div_p;
	wire dec_div_cancel;
	wire [31:0] exu_div_result;
	wire exu_div_wren;
	wire dec_i0_decode_d;
	wire [31:1] pred_correct_npc_x;
	wire [6:0] dec_tlu_br0_r_pkt;
	wire [55:0] exu_mp_pkt;
	wire [pt[2236-:8] - 1:0] exu_mp_eghr;
	wire [pt[2236-:8] - 1:0] exu_mp_fghr;
	wire [pt[2172-:9]:pt[2163-:6]] exu_mp_index;
	wire [pt[2139-:9] - 1:0] exu_mp_btag;
	wire [pt[2236-:8] - 1:0] exu_i0_br_fghr_r;
	wire [1:0] exu_i0_br_hist_r;
	wire exu_i0_br_error_r;
	wire exu_i0_br_start_error_r;
	wire exu_i0_br_valid_r;
	wire exu_i0_br_mp_r;
	wire exu_i0_br_middle_r;
	wire exu_i0_br_way_r;
	wire [pt[2172-:9]:pt[2163-:6]] exu_i0_br_index_r;
	wire dma_dccm_req;
	wire dma_iccm_req;
	wire [2:0] dma_mem_tag;
	wire [31:0] dma_mem_addr;
	wire [2:0] dma_mem_sz;
	wire dma_mem_write;
	wire [63:0] dma_mem_wdata;
	wire dccm_dma_rvalid;
	wire dccm_dma_ecc_error;
	wire [2:0] dccm_dma_rtag;
	wire [63:0] dccm_dma_rdata;
	wire iccm_dma_rvalid;
	wire iccm_dma_ecc_error;
	wire [2:0] iccm_dma_rtag;
	wire [63:0] iccm_dma_rdata;
	wire dma_dccm_stall_any;
	wire dma_iccm_stall_any;
	wire dccm_ready;
	wire iccm_ready;
	wire dma_pmu_dccm_read;
	wire dma_pmu_dccm_write;
	wire dma_pmu_any_read;
	wire dma_pmu_any_write;
	wire ifu_i0_icaf;
	wire [1:0] ifu_i0_icaf_type;
	wire ifu_i0_icaf_second;
	wire ifu_i0_dbecc;
	wire iccm_dma_sb_error;
	wire [50:0] i0_brp;
	wire [pt[2172-:9]:pt[2163-:6]] ifu_i0_bp_index;
	wire [pt[2236-:8] - 1:0] ifu_i0_bp_fghr;
	wire [pt[2139-:9] - 1:0] ifu_i0_bp_btag;
	wire [$clog2(pt[2061-:14]) - 1:0] ifu_i0_fa_index;
	wire [$clog2(pt[2061-:14]) - 1:0] dec_fa_error_index;
	wire [55:0] dec_i0_predict_p_d;
	wire [pt[2236-:8] - 1:0] i0_predict_fghr_d;
	wire [pt[2172-:9]:pt[2163-:6]] i0_predict_index_d;
	wire [pt[2139-:9] - 1:0] i0_predict_btag_d;
	wire picm_wren;
	wire picm_rden;
	wire picm_mken;
	wire [31:0] picm_rdaddr;
	wire [31:0] picm_wraddr;
	wire [31:0] picm_wr_data;
	wire [31:0] picm_rd_data;
	wire dec_tlu_external_ldfwd_disable;
	wire dec_tlu_bpred_disable;
	wire dec_tlu_wb_coalescing_disable;
	wire dec_tlu_sideeffect_posted_disable;
	wire [2:0] dec_tlu_dma_qos_prty;
	wire dec_tlu_misc_clk_override;
	wire dec_tlu_ifu_clk_override;
	wire dec_tlu_lsu_clk_override;
	wire dec_tlu_bus_clk_override;
	wire dec_tlu_pic_clk_override;
	wire dec_tlu_dccm_clk_override;
	wire dec_tlu_icm_clk_override;
	wire dec_tlu_picio_clk_override;
	assign dccm_clk_override = dec_tlu_dccm_clk_override;
	assign icm_clk_override = dec_tlu_icm_clk_override;
	wire [31:0] dbg_cmd_addr;
	wire [31:0] dbg_cmd_wrdata;
	wire dbg_cmd_valid;
	wire dbg_cmd_write;
	wire [1:0] dbg_cmd_type;
	wire [1:0] dbg_cmd_size;
	wire dbg_halt_req;
	wire dbg_resume_req;
	wire dbg_core_rst_l;
	wire core_dbg_cmd_done;
	wire core_dbg_cmd_fail;
	wire [31:0] core_dbg_rddata;
	wire dma_dbg_cmd_done;
	wire dma_dbg_cmd_fail;
	wire [31:0] dma_dbg_rddata;
	wire dbg_dma_bubble;
	wire dma_dbg_ready;
	wire [31:0] dec_dbg_rddata;
	wire dec_dbg_cmd_done;
	wire dec_dbg_cmd_fail;
	wire dec_tlu_mpc_halted_only;
	wire dec_tlu_dbg_halted;
	wire dec_tlu_resume_ack;
	wire dec_tlu_debug_mode;
	wire dec_debug_wdata_rs1_d;
	wire dec_tlu_force_halt;
	wire [1:0] dec_data_en;
	wire [1:0] dec_ctl_en;
	wire exu_pmu_i0_br_misp;
	wire exu_pmu_i0_br_ataken;
	wire exu_pmu_i0_pc4;
	wire lsu_pmu_load_external_m;
	wire lsu_pmu_store_external_m;
	wire lsu_pmu_misaligned_m;
	wire lsu_pmu_bus_trxn;
	wire lsu_pmu_bus_misaligned;
	wire lsu_pmu_bus_error;
	wire lsu_pmu_bus_busy;
	wire ifu_pmu_fetch_stall;
	wire ifu_pmu_ic_miss;
	wire ifu_pmu_ic_hit;
	wire ifu_pmu_bus_error;
	wire ifu_pmu_bus_busy;
	wire ifu_pmu_bus_trxn;
	wire active_state;
	wire free_clk;
	wire active_clk;
	wire dec_pause_state_cg;
	wire lsu_nonblock_load_data_error;
	wire [15:0] ifu_i0_cinst;
	wire [31:2] dec_tlu_meihap;
	wire dec_extint_stall;
	wire [103:0] trace_rv_trace_pkt;
	wire lsu_fastint_stall_any;
	wire [7:0] pic_claimid;
	wire [3:0] pic_pl;
	wire [3:0] dec_tlu_meicurpl;
	wire [3:0] dec_tlu_meipt;
	wire mexintpend;
	wire mhwakeup;
	wire dma_active;
	wire pause_state;
	wire halt_state;
	wire dec_tlu_core_empty;
	assign pause_state = (dec_pause_state_cg & ~(dma_active | lsu_active)) & dec_tlu_core_empty;
	assign halt_state = o_cpu_halt_status & ~(dma_active | lsu_active);
	assign active_state = ((~(halt_state | pause_state) | dec_tlu_flush_lower_r) | dec_tlu_flush_lower_wb) | dec_tlu_misc_clk_override;
	rvoclkhdr free_cg2(
		.clk(clk),
		.en(1'b1),
		.l1clk(free_l2clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr active_cg2(
		.clk(clk),
		.en(active_state),
		.l1clk(active_l2clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr free_cg1(
		.clk(free_l2clk),
		.en(1'b1),
		.l1clk(free_clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr active_cg1(
		.clk(active_l2clk),
		.en(1'b1),
		.l1clk(active_clk),
		.scan_mode(scan_mode)
	);
	assign core_dbg_cmd_done = dma_dbg_cmd_done | dec_dbg_cmd_done;
	assign core_dbg_cmd_fail = dma_dbg_cmd_fail | dec_dbg_cmd_fail;
	assign core_dbg_rddata[31:0] = (dma_dbg_cmd_done ? dma_dbg_rddata[31:0] : dec_dbg_rddata[31:0]);
	eb1_dbg #(.pt(pt)) dbg(
		.rst_l(core_rst_l),
		.clk(free_l2clk),
		.clk_override(dec_tlu_misc_clk_override),
		.sb_axi_awready(sb_axi_awready_int),
		.sb_axi_wready(sb_axi_wready_int),
		.sb_axi_bvalid(sb_axi_bvalid_int),
		.sb_axi_bresp(sb_axi_bresp_int[1:0]),
		.sb_axi_arready(sb_axi_arready_int),
		.sb_axi_rvalid(sb_axi_rvalid_int),
		.sb_axi_rdata(sb_axi_rdata_int[63:0]),
		.sb_axi_rresp(sb_axi_rresp_int[1:0]),
		.dbg_cmd_addr(dbg_cmd_addr),
		.dbg_cmd_wrdata(dbg_cmd_wrdata),
		.dbg_cmd_valid(dbg_cmd_valid),
		.dbg_cmd_write(dbg_cmd_write),
		.dbg_cmd_type(dbg_cmd_type),
		.dbg_cmd_size(dbg_cmd_size),
		.dbg_core_rst_l(dbg_core_rst_l),
		.core_dbg_rddata(core_dbg_rddata),
		.core_dbg_cmd_done(core_dbg_cmd_done),
		.core_dbg_cmd_fail(core_dbg_cmd_fail),
		.dbg_dma_bubble(dbg_dma_bubble),
		.dma_dbg_ready(dma_dbg_ready),
		.dbg_halt_req(dbg_halt_req),
		.dbg_resume_req(dbg_resume_req),
		.dec_tlu_debug_mode(dec_tlu_debug_mode),
		.dec_tlu_dbg_halted(dec_tlu_dbg_halted),
		.dec_tlu_mpc_halted_only(dec_tlu_mpc_halted_only),
		.dec_tlu_resume_ack(dec_tlu_resume_ack),
		.dmi_reg_en(dmi_reg_en),
		.dmi_reg_addr(dmi_reg_addr),
		.dmi_reg_wr_en(dmi_reg_wr_en),
		.dmi_reg_wdata(dmi_reg_wdata),
		.dmi_reg_rdata(dmi_reg_rdata),
		.sb_axi_awvalid(sb_axi_awvalid),
		.sb_axi_awid(sb_axi_awid),
		.sb_axi_awaddr(sb_axi_awaddr),
		.sb_axi_awregion(sb_axi_awregion),
		.sb_axi_awlen(sb_axi_awlen),
		.sb_axi_awsize(sb_axi_awsize),
		.sb_axi_awburst(sb_axi_awburst),
		.sb_axi_awlock(sb_axi_awlock),
		.sb_axi_awcache(sb_axi_awcache),
		.sb_axi_awprot(sb_axi_awprot),
		.sb_axi_awqos(sb_axi_awqos),
		.sb_axi_wvalid(sb_axi_wvalid),
		.sb_axi_wdata(sb_axi_wdata),
		.sb_axi_wstrb(sb_axi_wstrb),
		.sb_axi_wlast(sb_axi_wlast),
		.sb_axi_bready(sb_axi_bready),
		.sb_axi_arvalid(sb_axi_arvalid),
		.sb_axi_arid(sb_axi_arid),
		.sb_axi_araddr(sb_axi_araddr),
		.sb_axi_arregion(sb_axi_arregion),
		.sb_axi_arlen(sb_axi_arlen),
		.sb_axi_arsize(sb_axi_arsize),
		.sb_axi_arburst(sb_axi_arburst),
		.sb_axi_arlock(sb_axi_arlock),
		.sb_axi_arcache(sb_axi_arcache),
		.sb_axi_arprot(sb_axi_arprot),
		.sb_axi_arqos(sb_axi_arqos),
		.sb_axi_rready(sb_axi_rready),
		.dbg_bus_clk_en(dbg_bus_clk_en),
		.dbg_rst_l(dbg_rst_l),
		.scan_mode(scan_mode)
	);
	assign core_rst_l = rst_l & (dbg_core_rst_l | scan_mode);
	eb1_ifu #(.pt(pt)) ifu(
		.clk(active_l2clk),
		.rst_l(core_rst_l),
		.dec_tlu_flush_err_wb(dec_tlu_flush_err_r),
		.dec_tlu_flush_noredir_wb(dec_tlu_flush_noredir_r),
		.dec_tlu_fence_i_wb(dec_tlu_fence_i_r),
		.dec_tlu_flush_leak_one_wb(dec_tlu_flush_leak_one_r),
		.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_r),
		.ifu_axi_arready(ifu_axi_arready_int),
		.ifu_axi_rvalid(ifu_axi_rvalid_int),
		.ifu_axi_rid(ifu_axi_rid_int[pt[826-:8] - 1:0]),
		.ifu_axi_rdata(ifu_axi_rdata_int[63:0]),
		.ifu_axi_rresp(ifu_axi_rresp_int[1:0]),
		.exu_flush_final(exu_flush_final),
		.free_l2clk(free_l2clk),
		.active_clk(active_clk),
		.dec_i0_decode_d(dec_i0_decode_d),
		.dec_tlu_i0_commit_cmt(dec_tlu_i0_commit_cmt),
		.exu_flush_path_final(exu_flush_path_final),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.dec_tlu_bpred_disable(dec_tlu_bpred_disable),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.ifu_axi_awvalid(ifu_axi_awvalid),
		.ifu_axi_awid(ifu_axi_awid),
		.ifu_axi_awaddr(ifu_axi_awaddr),
		.ifu_axi_awregion(ifu_axi_awregion),
		.ifu_axi_awlen(ifu_axi_awlen),
		.ifu_axi_awsize(ifu_axi_awsize),
		.ifu_axi_awburst(ifu_axi_awburst),
		.ifu_axi_awlock(ifu_axi_awlock),
		.ifu_axi_awcache(ifu_axi_awcache),
		.ifu_axi_awprot(ifu_axi_awprot),
		.ifu_axi_awqos(ifu_axi_awqos),
		.ifu_axi_wvalid(ifu_axi_wvalid),
		.ifu_axi_wdata(ifu_axi_wdata),
		.ifu_axi_wstrb(ifu_axi_wstrb),
		.ifu_axi_wlast(ifu_axi_wlast),
		.ifu_axi_bready(ifu_axi_bready),
		.ifu_axi_arvalid(ifu_axi_arvalid),
		.ifu_axi_arid(ifu_axi_arid),
		.ifu_axi_araddr(ifu_axi_araddr),
		.ifu_axi_arregion(ifu_axi_arregion),
		.ifu_axi_arlen(ifu_axi_arlen),
		.ifu_axi_arsize(ifu_axi_arsize),
		.ifu_axi_arburst(ifu_axi_arburst),
		.ifu_axi_arlock(ifu_axi_arlock),
		.ifu_axi_arcache(ifu_axi_arcache),
		.ifu_axi_arprot(ifu_axi_arprot),
		.ifu_axi_arqos(ifu_axi_arqos),
		.ifu_axi_rready(ifu_axi_rready),
		.ifu_bus_clk_en(ifu_bus_clk_en),
		.dma_iccm_req(dma_iccm_req),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_sz(dma_mem_sz),
		.dma_mem_write(dma_mem_write),
		.dma_mem_wdata(dma_mem_wdata),
		.dma_mem_tag(dma_mem_tag),
		.dma_iccm_stall_any(dma_iccm_stall_any),
		.iccm_dma_ecc_error(iccm_dma_ecc_error),
		.iccm_dma_rvalid(iccm_dma_rvalid),
		.iccm_dma_rdata(iccm_dma_rdata),
		.iccm_dma_rtag(iccm_dma_rtag),
		.iccm_ready(iccm_ready),
		.ifu_pmu_instr_aligned(ifu_pmu_instr_aligned),
		.ifu_pmu_fetch_stall(ifu_pmu_fetch_stall),
		.ifu_ic_error_start(ifu_ic_error_start),
		.ic_rw_addr(ic_rw_addr),
		.ic_wr_en(ic_wr_en),
		.ic_rd_en(ic_rd_en),
		.ic_wr_data(ic_wr_data),
		.ic_rd_data(ic_rd_data),
		.ic_debug_rd_data(ic_debug_rd_data),
		.ictag_debug_rd_data(ictag_debug_rd_data),
		.ic_debug_wr_data(ic_debug_wr_data),
		.ifu_ic_debug_rd_data(ifu_ic_debug_rd_data),
		.ic_eccerr(ic_eccerr),
		.ic_parerr(ic_parerr),
		.ic_premux_data(ic_premux_data),
		.ic_sel_premux_data(ic_sel_premux_data),
		.ic_debug_addr(ic_debug_addr),
		.ic_debug_rd_en(ic_debug_rd_en),
		.ic_debug_wr_en(ic_debug_wr_en),
		.ic_debug_tag_array(ic_debug_tag_array),
		.ic_debug_way(ic_debug_way),
		.ic_tag_valid(ic_tag_valid),
		.ic_rd_hit(ic_rd_hit),
		.ic_tag_perr(ic_tag_perr),
		.iccm_rw_addr(iccm_rw_addr),
		.iccm_wren(iccm_wren),
		.iccm_rden(iccm_rden),
		.iccm_wr_data(iccm_wr_data),
		.iccm_wr_size(iccm_wr_size),
		.iccm_rd_data(iccm_rd_data),
		.iccm_rd_data_ecc(iccm_rd_data_ecc),
		.ifu_iccm_rd_ecc_single_err(ifu_iccm_rd_ecc_single_err),
		.ifu_pmu_ic_miss(ifu_pmu_ic_miss),
		.ifu_pmu_ic_hit(ifu_pmu_ic_hit),
		.ifu_pmu_bus_error(ifu_pmu_bus_error),
		.ifu_pmu_bus_busy(ifu_pmu_bus_busy),
		.ifu_pmu_bus_trxn(ifu_pmu_bus_trxn),
		.ifu_i0_icaf(ifu_i0_icaf),
		.ifu_i0_icaf_type(ifu_i0_icaf_type),
		.ifu_i0_valid(ifu_i0_valid),
		.ifu_i0_icaf_second(ifu_i0_icaf_second),
		.ifu_i0_dbecc(ifu_i0_dbecc),
		.iccm_dma_sb_error(iccm_dma_sb_error),
		.ifu_i0_instr(ifu_i0_instr),
		.ifu_i0_pc(ifu_i0_pc),
		.ifu_i0_pc4(ifu_i0_pc4),
		.ifu_miss_state_idle(ifu_miss_state_idle),
		.i0_brp(i0_brp),
		.ifu_i0_bp_index(ifu_i0_bp_index),
		.ifu_i0_bp_fghr(ifu_i0_bp_fghr),
		.ifu_i0_bp_btag(ifu_i0_bp_btag),
		.ifu_i0_fa_index(ifu_i0_fa_index),
		.exu_mp_pkt(exu_mp_pkt),
		.exu_mp_eghr(exu_mp_eghr),
		.exu_mp_fghr(exu_mp_fghr),
		.exu_mp_index(exu_mp_index),
		.exu_mp_btag(exu_mp_btag),
		.dec_tlu_br0_r_pkt(dec_tlu_br0_r_pkt),
		.exu_i0_br_fghr_r(exu_i0_br_fghr_r),
		.exu_i0_br_index_r(exu_i0_br_index_r),
		.dec_fa_error_index(dec_fa_error_index),
		.ifu_i0_cinst(ifu_i0_cinst),
		.dec_tlu_ic_diag_pkt(dec_tlu_ic_diag_pkt),
		.ifu_ic_debug_rd_data_valid(ifu_ic_debug_rd_data_valid),
		.iccm_buf_correct_ecc(iccm_buf_correct_ecc),
		.iccm_correction_state(iccm_correction_state),
		.scan_mode(scan_mode)
	);
	eb1_dec #(.pt(pt)) dec(
		.clk(active_l2clk),
		.dbg_cmd_wrdata(dbg_cmd_wrdata[1:0]),
		.rst_l(core_rst_l),
		.i_cpu_halt_req(i_cpu_halt_req),
		.i_cpu_run_req(i_cpu_run_req),
		.active_clk(active_clk),
		.free_clk(free_clk),
		.free_l2clk(free_l2clk),
		.lsu_fastint_stall_any(lsu_fastint_stall_any),
		.dec_extint_stall(dec_extint_stall),
		.dec_i0_decode_d(dec_i0_decode_d),
		.dec_pause_state_cg(dec_pause_state_cg),
		.dec_tlu_core_empty(dec_tlu_core_empty),
		.rst_vec(rst_vec),
		.nmi_int(nmi_int),
		.nmi_vec(nmi_vec),
		.o_cpu_halt_status(o_cpu_halt_status),
		.o_cpu_halt_ack(o_cpu_halt_ack),
		.o_cpu_run_ack(o_cpu_run_ack),
		.o_debug_mode_status(o_debug_mode_status),
		.core_id(core_id),
		.mpc_debug_halt_req(mpc_debug_halt_req),
		.mpc_debug_run_req(mpc_debug_run_req),
		.mpc_reset_run_req(mpc_reset_run_req),
		.mpc_debug_halt_ack(mpc_debug_halt_ack),
		.mpc_debug_run_ack(mpc_debug_run_ack),
		.debug_brkpt_status(debug_brkpt_status),
		.exu_pmu_i0_br_misp(exu_pmu_i0_br_misp),
		.exu_pmu_i0_br_ataken(exu_pmu_i0_br_ataken),
		.exu_pmu_i0_pc4(exu_pmu_i0_pc4),
		.lsu_nonblock_load_valid_m(lsu_nonblock_load_valid_m),
		.lsu_nonblock_load_tag_m(lsu_nonblock_load_tag_m),
		.lsu_nonblock_load_inv_r(lsu_nonblock_load_inv_r),
		.lsu_nonblock_load_inv_tag_r(lsu_nonblock_load_inv_tag_r),
		.lsu_nonblock_load_data_valid(lsu_nonblock_load_data_valid),
		.lsu_nonblock_load_data_error(lsu_nonblock_load_data_error),
		.lsu_nonblock_load_data_tag(lsu_nonblock_load_data_tag),
		.lsu_nonblock_load_data(lsu_nonblock_load_data),
		.lsu_pmu_bus_trxn(lsu_pmu_bus_trxn),
		.lsu_pmu_bus_misaligned(lsu_pmu_bus_misaligned),
		.lsu_pmu_bus_error(lsu_pmu_bus_error),
		.lsu_pmu_bus_busy(lsu_pmu_bus_busy),
		.lsu_pmu_misaligned_m(lsu_pmu_misaligned_m),
		.lsu_pmu_load_external_m(lsu_pmu_load_external_m),
		.lsu_pmu_store_external_m(lsu_pmu_store_external_m),
		.dma_pmu_dccm_read(dma_pmu_dccm_read),
		.dma_pmu_dccm_write(dma_pmu_dccm_write),
		.dma_pmu_any_read(dma_pmu_any_read),
		.dma_pmu_any_write(dma_pmu_any_write),
		.lsu_fir_addr(lsu_fir_addr),
		.lsu_fir_error(lsu_fir_error),
		.ifu_pmu_instr_aligned(ifu_pmu_instr_aligned),
		.ifu_pmu_fetch_stall(ifu_pmu_fetch_stall),
		.ifu_pmu_ic_miss(ifu_pmu_ic_miss),
		.ifu_pmu_ic_hit(ifu_pmu_ic_hit),
		.ifu_pmu_bus_error(ifu_pmu_bus_error),
		.ifu_pmu_bus_busy(ifu_pmu_bus_busy),
		.ifu_pmu_bus_trxn(ifu_pmu_bus_trxn),
		.ifu_ic_error_start(ifu_ic_error_start),
		.ifu_iccm_rd_ecc_single_err(ifu_iccm_rd_ecc_single_err),
		.lsu_trigger_match_m(lsu_trigger_match_m),
		.dbg_cmd_valid(dbg_cmd_valid),
		.dbg_cmd_write(dbg_cmd_write),
		.dbg_cmd_type(dbg_cmd_type),
		.dbg_cmd_addr(dbg_cmd_addr),
		.ifu_i0_icaf(ifu_i0_icaf),
		.ifu_i0_icaf_type(ifu_i0_icaf_type),
		.ifu_i0_icaf_second(ifu_i0_icaf_second),
		.ifu_i0_dbecc(ifu_i0_dbecc),
		.lsu_idle_any(lsu_idle_any),
		.i0_brp(i0_brp),
		.ifu_i0_bp_index(ifu_i0_bp_index),
		.ifu_i0_bp_fghr(ifu_i0_bp_fghr),
		.ifu_i0_bp_btag(ifu_i0_bp_btag),
		.ifu_i0_fa_index(ifu_i0_fa_index),
		.lsu_error_pkt_r(lsu_error_pkt_r),
		.lsu_single_ecc_error_incr(lsu_single_ecc_error_incr),
		.lsu_imprecise_error_load_any(lsu_imprecise_error_load_any),
		.lsu_imprecise_error_store_any(lsu_imprecise_error_store_any),
		.lsu_imprecise_error_addr_any(lsu_imprecise_error_addr_any),
		.exu_div_result(exu_div_result),
		.exu_div_wren(exu_div_wren),
		.exu_csr_rs1_x(exu_csr_rs1_x),
		.lsu_result_m(lsu_result_m),
		.lsu_result_corr_r(lsu_result_corr_r),
		.lsu_load_stall_any(lsu_load_stall_any),
		.lsu_store_stall_any(lsu_store_stall_any),
		.dma_dccm_stall_any(dma_dccm_stall_any),
		.dma_iccm_stall_any(dma_iccm_stall_any),
		.iccm_dma_sb_error(iccm_dma_sb_error),
		.exu_flush_final(exu_flush_final),
		.exu_npc_r(exu_npc_r),
		.exu_i0_result_x(exu_i0_result_x),
		.ifu_i0_valid(ifu_i0_valid),
		.ifu_i0_instr(ifu_i0_instr),
		.ifu_i0_pc(ifu_i0_pc),
		.ifu_i0_pc4(ifu_i0_pc4),
		.exu_i0_pc_x(exu_i0_pc_x),
		.mexintpend(mexintpend),
		.timer_int(timer_int),
		.soft_int(soft_int),
		.pic_claimid(pic_claimid),
		.pic_pl(pic_pl),
		.mhwakeup(mhwakeup),
		.dec_tlu_meicurpl(dec_tlu_meicurpl),
		.dec_tlu_meipt(dec_tlu_meipt),
		.ifu_ic_debug_rd_data(ifu_ic_debug_rd_data),
		.ifu_ic_debug_rd_data_valid(ifu_ic_debug_rd_data_valid),
		.dec_tlu_ic_diag_pkt(dec_tlu_ic_diag_pkt),
		.dbg_halt_req(dbg_halt_req),
		.dbg_resume_req(dbg_resume_req),
		.ifu_miss_state_idle(ifu_miss_state_idle),
		.dec_tlu_dbg_halted(dec_tlu_dbg_halted),
		.dec_tlu_debug_mode(dec_tlu_debug_mode),
		.dec_tlu_resume_ack(dec_tlu_resume_ack),
		.dec_tlu_flush_noredir_r(dec_tlu_flush_noredir_r),
		.dec_tlu_mpc_halted_only(dec_tlu_mpc_halted_only),
		.dec_tlu_flush_leak_one_r(dec_tlu_flush_leak_one_r),
		.dec_tlu_flush_err_r(dec_tlu_flush_err_r),
		.dec_tlu_meihap(dec_tlu_meihap),
		.dec_debug_wdata_rs1_d(dec_debug_wdata_rs1_d),
		.dec_dbg_rddata(dec_dbg_rddata),
		.dec_dbg_cmd_done(dec_dbg_cmd_done),
		.dec_dbg_cmd_fail(dec_dbg_cmd_fail),
		.trigger_pkt_any(trigger_pkt_any),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.exu_i0_br_hist_r(exu_i0_br_hist_r),
		.exu_i0_br_error_r(exu_i0_br_error_r),
		.exu_i0_br_start_error_r(exu_i0_br_start_error_r),
		.exu_i0_br_valid_r(exu_i0_br_valid_r),
		.exu_i0_br_mp_r(exu_i0_br_mp_r),
		.exu_i0_br_middle_r(exu_i0_br_middle_r),
		.exu_i0_br_way_r(exu_i0_br_way_r),
		.dec_i0_rs1_en_d(dec_i0_rs1_en_d),
		.dec_i0_rs2_en_d(dec_i0_rs2_en_d),
		.gpr_i0_rs1_d(gpr_i0_rs1_d),
		.gpr_i0_rs2_d(gpr_i0_rs2_d),
		.dec_i0_immed_d(dec_i0_immed_d),
		.dec_i0_br_immed_d(dec_i0_br_immed_d),
		.i0_ap(i0_ap),
		.dec_i0_alu_decode_d(dec_i0_alu_decode_d),
		.dec_i0_branch_d(dec_i0_branch_d),
		.dec_i0_select_pc_d(dec_i0_select_pc_d),
		.dec_i0_pc_d(dec_i0_pc_d),
		.dec_i0_rs1_bypass_en_d(dec_i0_rs1_bypass_en_d),
		.dec_i0_rs2_bypass_en_d(dec_i0_rs2_bypass_en_d),
		.dec_i0_result_r(dec_i0_result_r),
		.lsu_p(lsu_p),
		.dec_qual_lsu_d(dec_qual_lsu_d),
		.mul_p(mul_p),
		.div_p(div_p),
		.dec_div_cancel(dec_div_cancel),
		.dec_lsu_offset_d(dec_lsu_offset_d),
		.dec_csr_ren_d(dec_csr_ren_d),
		.dec_csr_rddata_d(dec_csr_rddata_d),
		.dec_tlu_flush_lower_r(dec_tlu_flush_lower_r),
		.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_wb),
		.dec_tlu_flush_path_r(dec_tlu_flush_path_r),
		.dec_tlu_i0_kill_writeb_r(dec_tlu_i0_kill_writeb_r),
		.dec_tlu_fence_i_r(dec_tlu_fence_i_r),
		.pred_correct_npc_x(pred_correct_npc_x),
		.dec_tlu_br0_r_pkt(dec_tlu_br0_r_pkt),
		.dec_tlu_perfcnt0(dec_tlu_perfcnt0),
		.dec_tlu_perfcnt1(dec_tlu_perfcnt1),
		.dec_tlu_perfcnt2(dec_tlu_perfcnt2),
		.dec_tlu_perfcnt3(dec_tlu_perfcnt3),
		.dec_i0_predict_p_d(dec_i0_predict_p_d),
		.i0_predict_fghr_d(i0_predict_fghr_d),
		.i0_predict_index_d(i0_predict_index_d),
		.i0_predict_btag_d(i0_predict_btag_d),
		.dec_fa_error_index(dec_fa_error_index),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.dec_data_en(dec_data_en),
		.dec_ctl_en(dec_ctl_en),
		.ifu_i0_cinst(ifu_i0_cinst),
		.trace_rv_trace_pkt(trace_rv_trace_pkt),
		.dec_tlu_external_ldfwd_disable(dec_tlu_external_ldfwd_disable),
		.dec_tlu_sideeffect_posted_disable(dec_tlu_sideeffect_posted_disable),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.dec_tlu_bpred_disable(dec_tlu_bpred_disable),
		.dec_tlu_wb_coalescing_disable(dec_tlu_wb_coalescing_disable),
		.dec_tlu_dma_qos_prty(dec_tlu_dma_qos_prty),
		.dec_tlu_misc_clk_override(dec_tlu_misc_clk_override),
		.dec_tlu_ifu_clk_override(dec_tlu_ifu_clk_override),
		.dec_tlu_lsu_clk_override(dec_tlu_lsu_clk_override),
		.dec_tlu_bus_clk_override(dec_tlu_bus_clk_override),
		.dec_tlu_pic_clk_override(dec_tlu_pic_clk_override),
		.dec_tlu_picio_clk_override(dec_tlu_picio_clk_override),
		.dec_tlu_dccm_clk_override(dec_tlu_dccm_clk_override),
		.dec_tlu_icm_clk_override(dec_tlu_icm_clk_override),
		.dec_tlu_i0_commit_cmt(dec_tlu_i0_commit_cmt),
		.scan_mode(scan_mode)
	);
	eb1_exu #(.pt(pt)) exu(
		.clk(active_l2clk),
		.rst_l(core_rst_l),
		.scan_mode(scan_mode),
		.dec_data_en(dec_data_en),
		.dec_ctl_en(dec_ctl_en),
		.dbg_cmd_wrdata(dbg_cmd_wrdata),
		.i0_ap(i0_ap),
		.dec_debug_wdata_rs1_d(dec_debug_wdata_rs1_d),
		.dec_i0_predict_p_d(dec_i0_predict_p_d),
		.i0_predict_fghr_d(i0_predict_fghr_d),
		.i0_predict_index_d(i0_predict_index_d),
		.i0_predict_btag_d(i0_predict_btag_d),
		.lsu_result_m(lsu_result_m),
		.lsu_nonblock_load_data(lsu_nonblock_load_data),
		.dec_i0_rs1_en_d(dec_i0_rs1_en_d),
		.dec_i0_rs2_en_d(dec_i0_rs2_en_d),
		.gpr_i0_rs1_d(gpr_i0_rs1_d),
		.gpr_i0_rs2_d(gpr_i0_rs2_d),
		.dec_i0_immed_d(dec_i0_immed_d),
		.dec_i0_result_r(dec_i0_result_r),
		.dec_i0_br_immed_d(dec_i0_br_immed_d),
		.dec_i0_alu_decode_d(dec_i0_alu_decode_d),
		.dec_i0_branch_d(dec_i0_branch_d),
		.dec_i0_select_pc_d(dec_i0_select_pc_d),
		.dec_i0_pc_d(dec_i0_pc_d),
		.dec_i0_rs1_bypass_en_d(dec_i0_rs1_bypass_en_d),
		.dec_i0_rs2_bypass_en_d(dec_i0_rs2_bypass_en_d),
		.dec_csr_ren_d(dec_csr_ren_d),
		.dec_csr_rddata_d(dec_csr_rddata_d),
		.dec_qual_lsu_d(dec_qual_lsu_d),
		.mul_p(mul_p),
		.div_p(div_p),
		.dec_div_cancel(dec_div_cancel),
		.pred_correct_npc_x(pred_correct_npc_x),
		.dec_tlu_flush_lower_r(dec_tlu_flush_lower_r),
		.dec_tlu_flush_path_r(dec_tlu_flush_path_r),
		.dec_extint_stall(dec_extint_stall),
		.dec_tlu_meihap(dec_tlu_meihap),
		.exu_lsu_rs1_d(exu_lsu_rs1_d),
		.exu_lsu_rs2_d(exu_lsu_rs2_d),
		.exu_flush_final(exu_flush_final),
		.exu_flush_path_final(exu_flush_path_final),
		.exu_i0_result_x(exu_i0_result_x),
		.exu_i0_pc_x(exu_i0_pc_x),
		.exu_csr_rs1_x(exu_csr_rs1_x),
		.exu_npc_r(exu_npc_r),
		.exu_i0_br_hist_r(exu_i0_br_hist_r),
		.exu_i0_br_error_r(exu_i0_br_error_r),
		.exu_i0_br_start_error_r(exu_i0_br_start_error_r),
		.exu_i0_br_index_r(exu_i0_br_index_r),
		.exu_i0_br_valid_r(exu_i0_br_valid_r),
		.exu_i0_br_mp_r(exu_i0_br_mp_r),
		.exu_i0_br_middle_r(exu_i0_br_middle_r),
		.exu_i0_br_fghr_r(exu_i0_br_fghr_r),
		.exu_i0_br_way_r(exu_i0_br_way_r),
		.exu_mp_pkt(exu_mp_pkt),
		.exu_mp_eghr(exu_mp_eghr),
		.exu_mp_fghr(exu_mp_fghr),
		.exu_mp_index(exu_mp_index),
		.exu_mp_btag(exu_mp_btag),
		.exu_pmu_i0_br_misp(exu_pmu_i0_br_misp),
		.exu_pmu_i0_br_ataken(exu_pmu_i0_br_ataken),
		.exu_pmu_i0_pc4(exu_pmu_i0_pc4),
		.exu_div_result(exu_div_result),
		.exu_div_wren(exu_div_wren)
	);
	eb1_lsu #(.pt(pt)) lsu(
		.clk(active_l2clk),
		.rst_l(core_rst_l),
		.clk_override(dec_tlu_lsu_clk_override),
		.dec_tlu_i0_kill_writeb_r(dec_tlu_i0_kill_writeb_r),
		.lsu_axi_awready(lsu_axi_awready_int),
		.lsu_axi_wready(lsu_axi_wready_int),
		.lsu_axi_bvalid(lsu_axi_bvalid_int),
		.lsu_axi_bid(lsu_axi_bid_int[pt[181-:8] - 1:0]),
		.lsu_axi_bresp(lsu_axi_bresp_int[1:0]),
		.lsu_axi_arready(lsu_axi_arready_int),
		.lsu_axi_rvalid(lsu_axi_rvalid_int),
		.lsu_axi_rid(lsu_axi_rid_int[pt[181-:8] - 1:0]),
		.lsu_axi_rdata(lsu_axi_rdata_int[63:0]),
		.lsu_axi_rresp(lsu_axi_rresp_int[1:0]),
		.lsu_axi_rlast(lsu_axi_rlast_int),
		.dec_tlu_flush_lower_r(dec_tlu_flush_lower_r),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.dec_tlu_external_ldfwd_disable(dec_tlu_external_ldfwd_disable),
		.dec_tlu_wb_coalescing_disable(dec_tlu_wb_coalescing_disable),
		.dec_tlu_sideeffect_posted_disable(dec_tlu_sideeffect_posted_disable),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.exu_lsu_rs1_d(exu_lsu_rs1_d),
		.exu_lsu_rs2_d(exu_lsu_rs2_d),
		.dec_lsu_offset_d(dec_lsu_offset_d),
		.lsu_p(lsu_p),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.lsu_result_m(lsu_result_m),
		.lsu_result_corr_r(lsu_result_corr_r),
		.lsu_load_stall_any(lsu_load_stall_any),
		.lsu_store_stall_any(lsu_store_stall_any),
		.lsu_fastint_stall_any(lsu_fastint_stall_any),
		.lsu_idle_any(lsu_idle_any),
		.lsu_active(lsu_active),
		.lsu_fir_addr(lsu_fir_addr),
		.lsu_fir_error(lsu_fir_error),
		.lsu_single_ecc_error_incr(lsu_single_ecc_error_incr),
		.lsu_error_pkt_r(lsu_error_pkt_r),
		.lsu_imprecise_error_load_any(lsu_imprecise_error_load_any),
		.lsu_imprecise_error_store_any(lsu_imprecise_error_store_any),
		.lsu_imprecise_error_addr_any(lsu_imprecise_error_addr_any),
		.lsu_nonblock_load_valid_m(lsu_nonblock_load_valid_m),
		.lsu_nonblock_load_tag_m(lsu_nonblock_load_tag_m),
		.lsu_nonblock_load_inv_r(lsu_nonblock_load_inv_r),
		.lsu_nonblock_load_inv_tag_r(lsu_nonblock_load_inv_tag_r),
		.lsu_nonblock_load_data_valid(lsu_nonblock_load_data_valid),
		.lsu_nonblock_load_data_error(lsu_nonblock_load_data_error),
		.lsu_nonblock_load_data_tag(lsu_nonblock_load_data_tag),
		.lsu_nonblock_load_data(lsu_nonblock_load_data),
		.lsu_pmu_load_external_m(lsu_pmu_load_external_m),
		.lsu_pmu_store_external_m(lsu_pmu_store_external_m),
		.lsu_pmu_misaligned_m(lsu_pmu_misaligned_m),
		.lsu_pmu_bus_trxn(lsu_pmu_bus_trxn),
		.lsu_pmu_bus_misaligned(lsu_pmu_bus_misaligned),
		.lsu_pmu_bus_error(lsu_pmu_bus_error),
		.lsu_pmu_bus_busy(lsu_pmu_bus_busy),
		.trigger_pkt_any(trigger_pkt_any),
		.lsu_trigger_match_m(lsu_trigger_match_m),
		.dccm_wren(dccm_wren),
		.dccm_rden(dccm_rden),
		.dccm_wr_addr_lo(dccm_wr_addr_lo),
		.dccm_wr_addr_hi(dccm_wr_addr_hi),
		.dccm_rd_addr_lo(dccm_rd_addr_lo),
		.dccm_rd_addr_hi(dccm_rd_addr_hi),
		.dccm_wr_data_lo(dccm_wr_data_lo),
		.dccm_wr_data_hi(dccm_wr_data_hi),
		.dccm_rd_data_lo(dccm_rd_data_lo),
		.dccm_rd_data_hi(dccm_rd_data_hi),
		.picm_wren(picm_wren),
		.picm_rden(picm_rden),
		.picm_mken(picm_mken),
		.picm_rdaddr(picm_rdaddr),
		.picm_wraddr(picm_wraddr),
		.picm_wr_data(picm_wr_data),
		.picm_rd_data(picm_rd_data),
		.lsu_axi_awvalid(lsu_axi_awvalid),
		.lsu_axi_awid(lsu_axi_awid),
		.lsu_axi_awaddr(lsu_axi_awaddr),
		.lsu_axi_awregion(lsu_axi_awregion),
		.lsu_axi_awlen(lsu_axi_awlen),
		.lsu_axi_awsize(lsu_axi_awsize),
		.lsu_axi_awburst(lsu_axi_awburst),
		.lsu_axi_awlock(lsu_axi_awlock),
		.lsu_axi_awcache(lsu_axi_awcache),
		.lsu_axi_awprot(lsu_axi_awprot),
		.lsu_axi_awqos(lsu_axi_awqos),
		.lsu_axi_wvalid(lsu_axi_wvalid),
		.lsu_axi_wdata(lsu_axi_wdata),
		.lsu_axi_wstrb(lsu_axi_wstrb),
		.lsu_axi_wlast(lsu_axi_wlast),
		.lsu_axi_bready(lsu_axi_bready),
		.lsu_axi_arvalid(lsu_axi_arvalid),
		.lsu_axi_arid(lsu_axi_arid),
		.lsu_axi_araddr(lsu_axi_araddr),
		.lsu_axi_arregion(lsu_axi_arregion),
		.lsu_axi_arlen(lsu_axi_arlen),
		.lsu_axi_arsize(lsu_axi_arsize),
		.lsu_axi_arburst(lsu_axi_arburst),
		.lsu_axi_arlock(lsu_axi_arlock),
		.lsu_axi_arcache(lsu_axi_arcache),
		.lsu_axi_arprot(lsu_axi_arprot),
		.lsu_axi_arqos(lsu_axi_arqos),
		.lsu_axi_rready(lsu_axi_rready),
		.lsu_bus_clk_en(lsu_bus_clk_en),
		.dma_dccm_req(dma_dccm_req),
		.dma_mem_tag(dma_mem_tag),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_sz(dma_mem_sz),
		.dma_mem_write(dma_mem_write),
		.dma_mem_wdata(dma_mem_wdata),
		.dccm_dma_rvalid(dccm_dma_rvalid),
		.dccm_dma_ecc_error(dccm_dma_ecc_error),
		.dccm_dma_rtag(dccm_dma_rtag),
		.dccm_dma_rdata(dccm_dma_rdata),
		.dccm_ready(dccm_ready),
		.scan_mode(scan_mode),
		.active_clk(active_clk)
	);
	eb1_pic_ctrl #(.pt(pt)) pic_ctrl_inst(
		.clk(free_l2clk),
		.clk_override(dec_tlu_pic_clk_override),
		.io_clk_override(dec_tlu_picio_clk_override),
		.picm_mken(picm_mken),
		.extintsrc_req({extintsrc_req[pt[56-:12]:1], 1'b0}),
		.pl(pic_pl[3:0]),
		.claimid(pic_claimid[7:0]),
		.meicurpl(dec_tlu_meicurpl[3:0]),
		.meipt(dec_tlu_meipt[3:0]),
		.rst_l(core_rst_l),
		.free_clk(free_clk),
		.picm_rdaddr(picm_rdaddr),
		.picm_wraddr(picm_wraddr),
		.picm_wr_data(picm_wr_data),
		.picm_wren(picm_wren),
		.picm_rden(picm_rden),
		.mexintpend(mexintpend),
		.picm_rd_data(picm_rd_data),
		.mhwakeup(mhwakeup),
		.scan_mode(scan_mode)
	);
	eb1_dma_ctrl #(.pt(pt)) dma_ctrl(
		.clk(free_l2clk),
		.rst_l(core_rst_l),
		.clk_override(dec_tlu_misc_clk_override),
		.dma_axi_awvalid(dma_axi_awvalid_int),
		.dma_axi_awid(dma_axi_awid_int[pt[1235-:8] - 1:0]),
		.dma_axi_awaddr(dma_axi_awaddr_int[31:0]),
		.dma_axi_awsize(dma_axi_awsize_int[2:0]),
		.dma_axi_wvalid(dma_axi_wvalid_int),
		.dma_axi_wdata(dma_axi_wdata_int[63:0]),
		.dma_axi_wstrb(dma_axi_wstrb_int[7:0]),
		.dma_axi_bready(dma_axi_bready_int),
		.dma_axi_arvalid(dma_axi_arvalid_int),
		.dma_axi_arid(dma_axi_arid_int[pt[1235-:8] - 1:0]),
		.dma_axi_araddr(dma_axi_araddr_int[31:0]),
		.dma_axi_arsize(dma_axi_arsize_int[2:0]),
		.dma_axi_rready(dma_axi_rready_int),
		.free_clk(free_clk),
		.dma_bus_clk_en(dma_bus_clk_en),
		.scan_mode(scan_mode),
		.dbg_cmd_addr(dbg_cmd_addr),
		.dbg_cmd_wrdata(dbg_cmd_wrdata),
		.dbg_cmd_valid(dbg_cmd_valid),
		.dbg_cmd_write(dbg_cmd_write),
		.dbg_cmd_type(dbg_cmd_type),
		.dbg_cmd_size(dbg_cmd_size),
		.dbg_dma_bubble(dbg_dma_bubble),
		.dma_dbg_ready(dma_dbg_ready),
		.dma_dbg_cmd_done(dma_dbg_cmd_done),
		.dma_dbg_cmd_fail(dma_dbg_cmd_fail),
		.dma_dbg_rddata(dma_dbg_rddata),
		.dma_dccm_req(dma_dccm_req),
		.dma_iccm_req(dma_iccm_req),
		.dma_mem_tag(dma_mem_tag),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_sz(dma_mem_sz),
		.dma_mem_write(dma_mem_write),
		.dma_mem_wdata(dma_mem_wdata),
		.dccm_dma_rvalid(dccm_dma_rvalid),
		.dccm_dma_ecc_error(dccm_dma_ecc_error),
		.dccm_dma_rtag(dccm_dma_rtag),
		.dccm_dma_rdata(dccm_dma_rdata),
		.iccm_dma_rvalid(iccm_dma_rvalid),
		.iccm_dma_ecc_error(iccm_dma_ecc_error),
		.iccm_dma_rtag(iccm_dma_rtag),
		.iccm_dma_rdata(iccm_dma_rdata),
		.dma_active(dma_active),
		.dma_dccm_stall_any(dma_dccm_stall_any),
		.dma_iccm_stall_any(dma_iccm_stall_any),
		.dccm_ready(dccm_ready),
		.iccm_ready(iccm_ready),
		.dec_tlu_dma_qos_prty(dec_tlu_dma_qos_prty),
		.dma_pmu_dccm_read(dma_pmu_dccm_read),
		.dma_pmu_dccm_write(dma_pmu_dccm_write),
		.dma_pmu_any_read(dma_pmu_any_read),
		.dma_pmu_any_write(dma_pmu_any_write),
		.dma_axi_awready(dma_axi_awready),
		.dma_axi_wready(dma_axi_wready),
		.dma_axi_bvalid(dma_axi_bvalid),
		.dma_axi_bresp(dma_axi_bresp),
		.dma_axi_bid(dma_axi_bid),
		.dma_axi_arready(dma_axi_arready),
		.dma_axi_rvalid(dma_axi_rvalid),
		.dma_axi_rid(dma_axi_rid),
		.dma_axi_rdata(dma_axi_rdata),
		.dma_axi_rresp(dma_axi_rresp),
		.dma_axi_rlast(dma_axi_rlast)
	);
	generate
		if (pt[2038] == 1) begin : Gen_AXI_To_AHB
			axi4_to_ahb #(
				.pt(pt),
				.TAG(pt[181-:8])
			) lsu_axi4_to_ahb(
				.clk(free_l2clk),
				.free_clk(free_clk),
				.rst_l(core_rst_l),
				.clk_override(dec_tlu_bus_clk_override),
				.bus_clk_en(lsu_bus_clk_en),
				.dec_tlu_force_halt(dec_tlu_force_halt),
				.axi_awvalid(lsu_axi_awvalid),
				.axi_awready(lsu_axi_awready_ahb),
				.axi_awid(lsu_axi_awid[pt[181-:8] - 1:0]),
				.axi_awaddr(lsu_axi_awaddr[31:0]),
				.axi_awsize(lsu_axi_awsize[2:0]),
				.axi_awprot(lsu_axi_awprot[2:0]),
				.axi_wvalid(lsu_axi_wvalid),
				.axi_wready(lsu_axi_wready_ahb),
				.axi_wdata(lsu_axi_wdata[63:0]),
				.axi_wstrb(lsu_axi_wstrb[7:0]),
				.axi_wlast(lsu_axi_wlast),
				.axi_bvalid(lsu_axi_bvalid_ahb),
				.axi_bready(lsu_axi_bready),
				.axi_bresp(lsu_axi_bresp_ahb[1:0]),
				.axi_bid(lsu_axi_bid_ahb[pt[181-:8] - 1:0]),
				.axi_arvalid(lsu_axi_arvalid),
				.axi_arready(lsu_axi_arready_ahb),
				.axi_arid(lsu_axi_arid[pt[181-:8] - 1:0]),
				.axi_araddr(lsu_axi_araddr[31:0]),
				.axi_arsize(lsu_axi_arsize[2:0]),
				.axi_arprot(lsu_axi_arprot[2:0]),
				.axi_rvalid(lsu_axi_rvalid_ahb),
				.axi_rready(lsu_axi_rready),
				.axi_rid(lsu_axi_rid_ahb[pt[181-:8] - 1:0]),
				.axi_rdata(lsu_axi_rdata_ahb[63:0]),
				.axi_rresp(lsu_axi_rresp_ahb[1:0]),
				.axi_rlast(lsu_axi_rlast_ahb),
				.ahb_haddr(lsu_haddr[31:0]),
				.ahb_hburst(lsu_hburst),
				.ahb_hmastlock(lsu_hmastlock),
				.ahb_hprot(lsu_hprot[3:0]),
				.ahb_hsize(lsu_hsize[2:0]),
				.ahb_htrans(lsu_htrans[1:0]),
				.ahb_hwrite(lsu_hwrite),
				.ahb_hwdata(lsu_hwdata[63:0]),
				.ahb_hrdata(lsu_hrdata[63:0]),
				.ahb_hready(lsu_hready),
				.ahb_hresp(lsu_hresp),
				.scan_mode(scan_mode)
			);
			axi4_to_ahb #(
				.pt(pt),
				.TAG(pt[826-:8])
			) ifu_axi4_to_ahb(
				.clk(free_l2clk),
				.free_clk(free_clk),
				.rst_l(core_rst_l),
				.clk_override(dec_tlu_bus_clk_override),
				.bus_clk_en(ifu_bus_clk_en),
				.dec_tlu_force_halt(dec_tlu_force_halt),
				.ahb_haddr(haddr[31:0]),
				.ahb_hburst(hburst),
				.ahb_hmastlock(hmastlock),
				.ahb_hprot(hprot[3:0]),
				.ahb_hsize(hsize[2:0]),
				.ahb_htrans(htrans[1:0]),
				.ahb_hwrite(hwrite),
				.ahb_hwdata(hwdata_nc[63:0]),
				.ahb_hrdata(hrdata[63:0]),
				.ahb_hready(hready),
				.ahb_hresp(hresp),
				.axi_awvalid(ifu_axi_awvalid),
				.axi_awready(ifu_axi_awready_ahb),
				.axi_awid(ifu_axi_awid[pt[826-:8] - 1:0]),
				.axi_awaddr(ifu_axi_awaddr[31:0]),
				.axi_awsize(ifu_axi_awsize[2:0]),
				.axi_awprot(ifu_axi_awprot[2:0]),
				.axi_wvalid(ifu_axi_wvalid),
				.axi_wready(ifu_axi_wready_ahb),
				.axi_wdata(ifu_axi_wdata[63:0]),
				.axi_wstrb(ifu_axi_wstrb[7:0]),
				.axi_wlast(ifu_axi_wlast),
				.axi_bvalid(ifu_axi_bvalid_ahb),
				.axi_bready(1'b1),
				.axi_bresp(ifu_axi_bresp_ahb[1:0]),
				.axi_bid(ifu_axi_bid_ahb[pt[826-:8] - 1:0]),
				.axi_arvalid(ifu_axi_arvalid),
				.axi_arready(ifu_axi_arready_ahb),
				.axi_arid(ifu_axi_arid[pt[826-:8] - 1:0]),
				.axi_araddr(ifu_axi_araddr[31:0]),
				.axi_arsize(ifu_axi_arsize[2:0]),
				.axi_arprot(ifu_axi_arprot[2:0]),
				.axi_rvalid(ifu_axi_rvalid_ahb),
				.axi_rready(ifu_axi_rready),
				.axi_rid(ifu_axi_rid_ahb[pt[826-:8] - 1:0]),
				.axi_rdata(ifu_axi_rdata_ahb[63:0]),
				.axi_rresp(ifu_axi_rresp_ahb[1:0]),
				.axi_rlast(ifu_axi_rlast_ahb),
				.scan_mode(scan_mode)
			);
			axi4_to_ahb #(
				.pt(pt),
				.TAG(pt[12-:8])
			) sb_axi4_to_ahb(
				.clk(free_l2clk),
				.free_clk(free_clk),
				.rst_l(dbg_rst_l),
				.clk_override(dec_tlu_bus_clk_override),
				.bus_clk_en(dbg_bus_clk_en),
				.dec_tlu_force_halt(1'b0),
				.axi_awvalid(sb_axi_awvalid),
				.axi_awready(sb_axi_awready_ahb),
				.axi_awid(sb_axi_awid[pt[12-:8] - 1:0]),
				.axi_awaddr(sb_axi_awaddr[31:0]),
				.axi_awsize(sb_axi_awsize[2:0]),
				.axi_awprot(sb_axi_awprot[2:0]),
				.axi_wvalid(sb_axi_wvalid),
				.axi_wready(sb_axi_wready_ahb),
				.axi_wdata(sb_axi_wdata[63:0]),
				.axi_wstrb(sb_axi_wstrb[7:0]),
				.axi_wlast(sb_axi_wlast),
				.axi_bvalid(sb_axi_bvalid_ahb),
				.axi_bready(sb_axi_bready),
				.axi_bresp(sb_axi_bresp_ahb[1:0]),
				.axi_bid(sb_axi_bid_ahb[pt[12-:8] - 1:0]),
				.axi_arvalid(sb_axi_arvalid),
				.axi_arready(sb_axi_arready_ahb),
				.axi_arid(sb_axi_arid[pt[12-:8] - 1:0]),
				.axi_araddr(sb_axi_araddr[31:0]),
				.axi_arsize(sb_axi_arsize[2:0]),
				.axi_arprot(sb_axi_arprot[2:0]),
				.axi_rvalid(sb_axi_rvalid_ahb),
				.axi_rready(sb_axi_rready),
				.axi_rid(sb_axi_rid_ahb[pt[12-:8] - 1:0]),
				.axi_rdata(sb_axi_rdata_ahb[63:0]),
				.axi_rresp(sb_axi_rresp_ahb[1:0]),
				.axi_rlast(sb_axi_rlast_ahb),
				.ahb_haddr(sb_haddr[31:0]),
				.ahb_hburst(sb_hburst),
				.ahb_hmastlock(sb_hmastlock),
				.ahb_hprot(sb_hprot[3:0]),
				.ahb_hsize(sb_hsize[2:0]),
				.ahb_htrans(sb_htrans[1:0]),
				.ahb_hwrite(sb_hwrite),
				.ahb_hwdata(sb_hwdata[63:0]),
				.ahb_hrdata(sb_hrdata[63:0]),
				.ahb_hready(sb_hready),
				.ahb_hresp(sb_hresp),
				.scan_mode(scan_mode)
			);
			ahb_to_axi4 #(
				.pt(pt),
				.TAG(pt[1235-:8])
			) dma_ahb_to_axi4(
				.clk(free_l2clk),
				.rst_l(core_rst_l),
				.clk_override(dec_tlu_bus_clk_override),
				.bus_clk_en(dma_bus_clk_en),
				.axi_awvalid(dma_axi_awvalid_ahb),
				.axi_awready(dma_axi_awready),
				.axi_awid(dma_axi_awid_ahb[pt[1235-:8] - 1:0]),
				.axi_awaddr(dma_axi_awaddr_ahb[31:0]),
				.axi_awsize(dma_axi_awsize_ahb[2:0]),
				.axi_awprot(dma_axi_awprot_ahb[2:0]),
				.axi_awlen(dma_axi_awlen_ahb[7:0]),
				.axi_awburst(dma_axi_awburst_ahb[1:0]),
				.axi_wvalid(dma_axi_wvalid_ahb),
				.axi_wready(dma_axi_wready),
				.axi_wdata(dma_axi_wdata_ahb[63:0]),
				.axi_wstrb(dma_axi_wstrb_ahb[7:0]),
				.axi_wlast(dma_axi_wlast_ahb),
				.axi_bvalid(dma_axi_bvalid),
				.axi_bready(dma_axi_bready_ahb),
				.axi_bresp(dma_axi_bresp[1:0]),
				.axi_bid(dma_axi_bid[pt[1235-:8] - 1:0]),
				.axi_arvalid(dma_axi_arvalid_ahb),
				.axi_arready(dma_axi_arready),
				.axi_arid(dma_axi_arid_ahb[pt[1235-:8] - 1:0]),
				.axi_araddr(dma_axi_araddr_ahb[31:0]),
				.axi_arsize(dma_axi_arsize_ahb[2:0]),
				.axi_arprot(dma_axi_arprot_ahb[2:0]),
				.axi_arlen(dma_axi_arlen_ahb[7:0]),
				.axi_arburst(dma_axi_arburst_ahb[1:0]),
				.axi_rvalid(dma_axi_rvalid),
				.axi_rready(dma_axi_rready_ahb),
				.axi_rid(dma_axi_rid[pt[1235-:8] - 1:0]),
				.axi_rdata(dma_axi_rdata[63:0]),
				.axi_rresp(dma_axi_rresp[1:0]),
				.ahb_haddr(dma_haddr[31:0]),
				.ahb_hburst(dma_hburst),
				.ahb_hmastlock(dma_hmastlock),
				.ahb_hprot(dma_hprot[3:0]),
				.ahb_hsize(dma_hsize[2:0]),
				.ahb_htrans(dma_htrans[1:0]),
				.ahb_hwrite(dma_hwrite),
				.ahb_hwdata(dma_hwdata[63:0]),
				.ahb_hrdata(dma_hrdata[63:0]),
				.ahb_hreadyout(dma_hreadyout),
				.ahb_hresp(dma_hresp),
				.ahb_hreadyin(dma_hreadyin),
				.ahb_hsel(dma_hsel),
				.scan_mode(scan_mode)
			);
		end
	endgenerate
	assign lsu_axi_awready_int = (pt[2038] ? lsu_axi_awready_ahb : lsu_axi_awready);
	assign lsu_axi_wready_int = (pt[2038] ? lsu_axi_wready_ahb : lsu_axi_wready);
	assign lsu_axi_bvalid_int = (pt[2038] ? lsu_axi_bvalid_ahb : lsu_axi_bvalid);
	assign lsu_axi_bready_int = (pt[2038] ? lsu_axi_bready_ahb : lsu_axi_bready);
	assign lsu_axi_bresp_int[1:0] = (pt[2038] ? lsu_axi_bresp_ahb[1:0] : lsu_axi_bresp[1:0]);
	assign lsu_axi_bid_int[pt[181-:8] - 1:0] = (pt[2038] ? lsu_axi_bid_ahb[pt[181-:8] - 1:0] : lsu_axi_bid[pt[181-:8] - 1:0]);
	assign lsu_axi_arready_int = (pt[2038] ? lsu_axi_arready_ahb : lsu_axi_arready);
	assign lsu_axi_rvalid_int = (pt[2038] ? lsu_axi_rvalid_ahb : lsu_axi_rvalid);
	assign lsu_axi_rid_int[pt[181-:8] - 1:0] = (pt[2038] ? lsu_axi_rid_ahb[pt[181-:8] - 1:0] : lsu_axi_rid[pt[181-:8] - 1:0]);
	assign lsu_axi_rdata_int[63:0] = (pt[2038] ? lsu_axi_rdata_ahb[63:0] : lsu_axi_rdata[63:0]);
	assign lsu_axi_rresp_int[1:0] = (pt[2038] ? lsu_axi_rresp_ahb[1:0] : lsu_axi_rresp[1:0]);
	assign lsu_axi_rlast_int = (pt[2038] ? lsu_axi_rlast_ahb : lsu_axi_rlast);
	assign ifu_axi_awready_int = (pt[2038] ? ifu_axi_awready_ahb : ifu_axi_awready);
	assign ifu_axi_wready_int = (pt[2038] ? ifu_axi_wready_ahb : ifu_axi_wready);
	assign ifu_axi_bvalid_int = (pt[2038] ? ifu_axi_bvalid_ahb : ifu_axi_bvalid);
	assign ifu_axi_bready_int = (pt[2038] ? ifu_axi_bready_ahb : ifu_axi_bready);
	assign ifu_axi_bresp_int[1:0] = (pt[2038] ? ifu_axi_bresp_ahb[1:0] : ifu_axi_bresp[1:0]);
	assign ifu_axi_bid_int[pt[826-:8] - 1:0] = (pt[2038] ? ifu_axi_bid_ahb[pt[826-:8] - 1:0] : ifu_axi_bid[pt[826-:8] - 1:0]);
	assign ifu_axi_arready_int = (pt[2038] ? ifu_axi_arready_ahb : ifu_axi_arready);
	assign ifu_axi_rvalid_int = (pt[2038] ? ifu_axi_rvalid_ahb : ifu_axi_rvalid);
	assign ifu_axi_rid_int[pt[826-:8] - 1:0] = (pt[2038] ? ifu_axi_rid_ahb[pt[826-:8] - 1:0] : ifu_axi_rid[pt[826-:8] - 1:0]);
	assign ifu_axi_rdata_int[63:0] = (pt[2038] ? ifu_axi_rdata_ahb[63:0] : ifu_axi_rdata[63:0]);
	assign ifu_axi_rresp_int[1:0] = (pt[2038] ? ifu_axi_rresp_ahb[1:0] : ifu_axi_rresp[1:0]);
	assign ifu_axi_rlast_int = (pt[2038] ? ifu_axi_rlast_ahb : ifu_axi_rlast);
	assign sb_axi_awready_int = (pt[2038] ? sb_axi_awready_ahb : sb_axi_awready);
	assign sb_axi_wready_int = (pt[2038] ? sb_axi_wready_ahb : sb_axi_wready);
	assign sb_axi_bvalid_int = (pt[2038] ? sb_axi_bvalid_ahb : sb_axi_bvalid);
	assign sb_axi_bready_int = (pt[2038] ? sb_axi_bready_ahb : sb_axi_bready);
	assign sb_axi_bresp_int[1:0] = (pt[2038] ? sb_axi_bresp_ahb[1:0] : sb_axi_bresp[1:0]);
	assign sb_axi_bid_int[pt[12-:8] - 1:0] = (pt[2038] ? sb_axi_bid_ahb[pt[12-:8] - 1:0] : sb_axi_bid[pt[12-:8] - 1:0]);
	assign sb_axi_arready_int = (pt[2038] ? sb_axi_arready_ahb : sb_axi_arready);
	assign sb_axi_rvalid_int = (pt[2038] ? sb_axi_rvalid_ahb : sb_axi_rvalid);
	assign sb_axi_rid_int[pt[12-:8] - 1:0] = (pt[2038] ? sb_axi_rid_ahb[pt[12-:8] - 1:0] : sb_axi_rid[pt[12-:8] - 1:0]);
	assign sb_axi_rdata_int[63:0] = (pt[2038] ? sb_axi_rdata_ahb[63:0] : sb_axi_rdata[63:0]);
	assign sb_axi_rresp_int[1:0] = (pt[2038] ? sb_axi_rresp_ahb[1:0] : sb_axi_rresp[1:0]);
	assign sb_axi_rlast_int = (pt[2038] ? sb_axi_rlast_ahb : sb_axi_rlast);
	assign dma_axi_awvalid_int = (pt[2038] ? dma_axi_awvalid_ahb : dma_axi_awvalid);
	assign dma_axi_awid_int[pt[1235-:8] - 1:0] = (pt[2038] ? dma_axi_awid_ahb[pt[1235-:8] - 1:0] : dma_axi_awid[pt[1235-:8] - 1:0]);
	assign dma_axi_awaddr_int[31:0] = (pt[2038] ? dma_axi_awaddr_ahb[31:0] : dma_axi_awaddr[31:0]);
	assign dma_axi_awsize_int[2:0] = (pt[2038] ? dma_axi_awsize_ahb[2:0] : dma_axi_awsize[2:0]);
	assign dma_axi_awprot_int[2:0] = (pt[2038] ? dma_axi_awprot_ahb[2:0] : dma_axi_awprot[2:0]);
	assign dma_axi_awlen_int[7:0] = (pt[2038] ? dma_axi_awlen_ahb[7:0] : dma_axi_awlen[7:0]);
	assign dma_axi_awburst_int[1:0] = (pt[2038] ? dma_axi_awburst_ahb[1:0] : dma_axi_awburst[1:0]);
	assign dma_axi_wvalid_int = (pt[2038] ? dma_axi_wvalid_ahb : dma_axi_wvalid);
	assign dma_axi_wdata_int[63:0] = (pt[2038] ? dma_axi_wdata_ahb[63:0] : dma_axi_wdata);
	assign dma_axi_wstrb_int[7:0] = (pt[2038] ? dma_axi_wstrb_ahb[7:0] : dma_axi_wstrb[7:0]);
	assign dma_axi_wlast_int = (pt[2038] ? dma_axi_wlast_ahb : dma_axi_wlast);
	assign dma_axi_bready_int = (pt[2038] ? dma_axi_bready_ahb : dma_axi_bready);
	assign dma_axi_arvalid_int = (pt[2038] ? dma_axi_arvalid_ahb : dma_axi_arvalid);
	assign dma_axi_arid_int[pt[1235-:8] - 1:0] = (pt[2038] ? dma_axi_arid_ahb[pt[1235-:8] - 1:0] : dma_axi_arid[pt[1235-:8] - 1:0]);
	assign dma_axi_araddr_int[31:0] = (pt[2038] ? dma_axi_araddr_ahb[31:0] : dma_axi_araddr[31:0]);
	assign dma_axi_arsize_int[2:0] = (pt[2038] ? dma_axi_arsize_ahb[2:0] : dma_axi_arsize[2:0]);
	assign dma_axi_arprot_int[2:0] = (pt[2038] ? dma_axi_arprot_ahb[2:0] : dma_axi_arprot[2:0]);
	assign dma_axi_arlen_int[7:0] = (pt[2038] ? dma_axi_arlen_ahb[7:0] : dma_axi_arlen[7:0]);
	assign dma_axi_arburst_int[1:0] = (pt[2038] ? dma_axi_arburst_ahb[1:0] : dma_axi_arburst[1:0]);
	assign dma_axi_rready_int = (pt[2038] ? dma_axi_rready_ahb : dma_axi_rready);
	assign trace_rv_i_insn_ip[31:0] = trace_rv_trace_pkt[102:71];
	assign trace_rv_i_address_ip[31:0] = trace_rv_trace_pkt[70:39];
	assign trace_rv_i_valid_ip = trace_rv_trace_pkt[103];
	assign trace_rv_i_exception_ip = trace_rv_trace_pkt[38];
	assign trace_rv_i_ecause_ip[4:0] = trace_rv_trace_pkt[37:33];
	assign trace_rv_i_interrupt_ip = trace_rv_trace_pkt[32];
	assign trace_rv_i_tval_ip[31:0] = trace_rv_trace_pkt[31:0];
endmodule
module dmi_wrapper (
	trst_n,
	tck,
	tms,
	tdi,
	tdo,
	tdoEnable,
	core_rst_n,
	core_clk,
	jtag_id,
	rd_data,
	reg_wr_data,
	reg_wr_addr,
	reg_en,
	reg_wr_en,
	dmi_hard_reset
);
	input trst_n;
	input tck;
	input tms;
	input tdi;
	output tdo;
	output tdoEnable;
	input core_rst_n;
	input core_clk;
	input [31:1] jtag_id;
	input [31:0] rd_data;
	output [31:0] reg_wr_data;
	output [6:0] reg_wr_addr;
	output reg_en;
	output reg_wr_en;
	output dmi_hard_reset;
	wire rd_en;
	wire wr_en;
	wire dmireset;
	rvjtag_tap i_jtag_tap(
		.trst(trst_n),
		.tck(tck),
		.tms(tms),
		.tdi(tdi),
		.tdo(tdo),
		.tdoEnable(tdoEnable),
		.wr_data(reg_wr_data),
		.wr_addr(reg_wr_addr),
		.rd_en(rd_en),
		.wr_en(wr_en),
		.rd_data(rd_data),
		.rd_status(2'b00),
		.idle(3'h0),
		.dmi_stat(2'b00),
		.version(4'h1),
		.jtag_id(jtag_id),
		.dmi_hard_reset(dmi_hard_reset),
		.dmi_reset(dmireset)
	);
	dmi_jtag_to_core_sync i_dmi_jtag_to_core_sync(
		.wr_en(wr_en),
		.rd_en(rd_en),
		.rst_n(core_rst_n),
		.clk(core_clk),
		.reg_en(reg_en),
		.reg_wr_en(reg_wr_en)
	);
endmodule
module eb1_uart_rx_prog (
	i_Clock,
	rst_ni,
	i_Rx_Serial,
	CLKS_PER_BIT,
	o_Rx_DV,
	o_Rx_Byte
);
	input i_Clock;
	input rst_ni;
	input i_Rx_Serial;
	input [15:0] CLKS_PER_BIT;
	output o_Rx_DV;
	output [7:0] o_Rx_Byte;
	parameter s_IDLE = 3'b000;
	parameter s_RX_START_BIT = 3'b001;
	parameter s_RX_DATA_BITS = 3'b010;
	parameter s_RX_STOP_BIT = 3'b011;
	parameter s_CLEANUP = 3'b100;
	reg r_Rx_Data_R;
	reg r_Rx_Data;
	reg [15:0] r_Clock_Count;
	reg [2:0] r_Bit_Index;
	reg [7:0] r_Rx_Byte;
	reg r_Rx_DV;
	reg [2:0] r_SM_Main;
	always @(posedge i_Clock)
		if (rst_ni == 1'b0) begin
			r_Rx_Data_R <= 1'b1;
			r_Rx_Data <= 1'b1;
		end
		else begin
			r_Rx_Data_R <= i_Rx_Serial;
			r_Rx_Data <= r_Rx_Data_R;
		end
	always @(posedge i_Clock or negedge rst_ni)
		if (rst_ni == 1'b0) begin
			r_SM_Main <= s_IDLE;
			r_Rx_DV <= 1'b0;
			r_Clock_Count <= 16'h0000;
			r_Bit_Index <= 3'b000;
			r_Rx_Byte <= 8'h00;
		end
		else
			case (r_SM_Main)
				s_IDLE: begin
					r_Rx_DV <= 1'b0;
					r_Clock_Count <= 0;
					r_Bit_Index <= 0;
					if (r_Rx_Data == 1'b0)
						r_SM_Main <= s_RX_START_BIT;
					else
						r_SM_Main <= s_IDLE;
				end
				s_RX_START_BIT:
					if (r_Clock_Count == ((CLKS_PER_BIT - 1) >> 1)) begin
						if (r_Rx_Data == 1'b0) begin
							r_Clock_Count <= 0;
							r_SM_Main <= s_RX_DATA_BITS;
						end
						else
							r_SM_Main <= s_IDLE;
					end
					else begin
						r_Clock_Count <= r_Clock_Count + 1;
						r_SM_Main <= s_RX_START_BIT;
					end
				s_RX_DATA_BITS:
					if (r_Clock_Count < (CLKS_PER_BIT - 1)) begin
						r_Clock_Count <= r_Clock_Count + 1;
						r_SM_Main <= s_RX_DATA_BITS;
					end
					else begin
						r_Clock_Count <= 0;
						r_Rx_Byte[r_Bit_Index] <= r_Rx_Data;
						if (r_Bit_Index < 7) begin
							r_Bit_Index <= r_Bit_Index + 1;
							r_SM_Main <= s_RX_DATA_BITS;
						end
						else begin
							r_Bit_Index <= 0;
							r_SM_Main <= s_RX_STOP_BIT;
						end
					end
				s_RX_STOP_BIT:
					if (r_Clock_Count < (CLKS_PER_BIT - 1)) begin
						r_Clock_Count <= r_Clock_Count + 1;
						r_SM_Main <= s_RX_STOP_BIT;
					end
					else begin
						r_Rx_DV <= 1'b1;
						r_Clock_Count <= 0;
						r_SM_Main <= s_CLEANUP;
					end
				s_CLEANUP: begin
					r_SM_Main <= s_IDLE;
					r_Rx_DV <= 1'b0;
				end
				default: r_SM_Main <= s_IDLE;
			endcase
	assign o_Rx_DV = r_Rx_DV;
	assign o_Rx_Byte = r_Rx_Byte;
endmodule
module eb1_iccm_controller (
	clk_i,
	rst_ni,
	rx_dv_i,
	rx_byte_i,
	we_o,
	addr_o,
	wdata_o,
	reset_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire rx_dv_i;
	input wire [7:0] rx_byte_i;
	output wire we_o;
	output wire [13:0] addr_o;
	output wire [31:0] wdata_o;
	output wire reset_o;
	reg [1:0] ctrl_fsm_cs;
	reg [1:0] ctrl_fsm_ns;
	wire [7:0] rx_byte_d;
	reg [7:0] rx_byte_q0;
	reg [7:0] rx_byte_q1;
	reg [7:0] rx_byte_q2;
	reg [7:0] rx_byte_q3;
	reg we_q;
	reg we_d;
	reg [13:0] addr_q;
	reg [13:0] addr_d;
	reg reset_q;
	reg reset_d;
	reg [1:0] byte_count;
	localparam [1:0] DONE = 3;
	localparam [1:0] LOAD = 1;
	localparam [1:0] PROG = 2;
	localparam [1:0] RESET = 0;
	always @(*) begin
		we_d = we_q;
		addr_d = addr_q;
		reset_d = reset_q;
		ctrl_fsm_ns = ctrl_fsm_cs;
		case (ctrl_fsm_cs)
			RESET: begin
				we_d = 1'b0;
				reset_d = 1'b0;
				if (rx_dv_i)
					ctrl_fsm_ns = LOAD;
				else
					ctrl_fsm_ns = RESET;
			end
			LOAD:
				if (((byte_count == 2'b11) && (rx_byte_q2 != 8'h0f)) && (rx_byte_d != 8'hff)) begin
					we_d = 1'b1;
					ctrl_fsm_ns = PROG;
				end
				else
					ctrl_fsm_ns = DONE;
			PROG: begin
				we_d = 1'b0;
				ctrl_fsm_ns = DONE;
			end
			DONE:
				if (wdata_o == 32'h00000fff) begin
					ctrl_fsm_ns = DONE;
					reset_d = 1'b1;
				end
				else if (rx_dv_i)
					ctrl_fsm_ns = LOAD;
				else
					ctrl_fsm_ns = DONE;
			default: ctrl_fsm_ns = RESET;
		endcase
	end
	assign rx_byte_d = rx_byte_i;
	assign we_o = we_q;
	assign addr_o = addr_q;
	assign wdata_o = {rx_byte_q0, rx_byte_q1, rx_byte_q2, rx_byte_q3};
	assign reset_o = reset_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			we_q <= 1'b0;
			addr_q <= 14'b00000000000000;
			rx_byte_q0 <= 8'b00000000;
			rx_byte_q1 <= 8'b00000000;
			rx_byte_q2 <= 8'b00000000;
			rx_byte_q3 <= 8'b00000000;
			reset_q <= 1'b0;
			byte_count <= 2'b00;
			ctrl_fsm_cs <= RESET;
		end
		else begin
			we_q <= we_d;
			if (ctrl_fsm_cs == LOAD) begin
				if (byte_count == 2'b00) begin
					rx_byte_q0 <= rx_byte_d;
					byte_count <= 2'b01;
				end
				else if (byte_count == 2'b01) begin
					rx_byte_q1 <= rx_byte_d;
					byte_count <= 2'b10;
				end
				else if (byte_count == 2'b10) begin
					rx_byte_q2 <= rx_byte_d;
					byte_count <= 2'b11;
				end
				else begin
					rx_byte_q3 <= rx_byte_d;
					byte_count <= 2'b00;
				end
				addr_q <= addr_d;
			end
			if (ctrl_fsm_cs == PROG)
				addr_q <= addr_d + 2'h2;
			reset_q <= reset_d;
			ctrl_fsm_cs <= ctrl_fsm_ns;
		end
endmodule
module eb1_mem (
`ifdef USE_POWER_PINS
	VPWR,
	VGND,
`endif
	clk,
	rst_l,
	dccm_clk_override,
	icm_clk_override,
	dec_tlu_core_ecc_disable,
	dccm_wren,
	dccm_rden,
	dccm_wr_addr_lo,
	dccm_wr_addr_hi,
	dccm_rd_addr_lo,
	dccm_rd_addr_hi,
	dccm_wr_data_lo,
	dccm_wr_data_hi,
	dccm_rd_data_lo,
	dccm_rd_data_hi,
	dccm_ext_in_pkt,
	iccm_ext_in_pkt,
	iccm_rw_addr,
	iccm_buf_correct_ecc,
	iccm_correction_state,
	iccm_wren,
	iccm_rden,
	iccm_wr_size,
	iccm_wr_data,
	iccm_rd_data,
	iccm_rd_data_ecc,
	ic_rw_addr,
	ic_tag_valid,
	ic_wr_en,
	ic_rd_en,
	ic_premux_data,
	ic_sel_premux_data,
	ic_data_ext_in_pkt,
	ic_tag_ext_in_pkt,
	ic_wr_data,
	ic_debug_wr_data,
	ic_debug_rd_data,
	ic_debug_addr,
	ic_debug_rd_en,
	ic_debug_wr_en,
	ic_debug_tag_array,
	ic_debug_way,
	ic_rd_data,
	ictag_debug_rd_data,
	ic_eccerr,
	ic_parerr,
	ic_rd_hit,
	ic_tag_perr,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
`ifdef USE_POWER_PINS
	inout wire VPWR;
	inout wire VGND;
`endif
	input wire clk;
	input wire rst_l;
	input wire dccm_clk_override;
	input wire icm_clk_override;
	input wire dec_tlu_core_ecc_disable;
	input wire dccm_wren;
	input wire dccm_rden;
	input wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	input wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	input wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	input wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	input wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	input wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	output wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	output wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	input wire [(pt[1342-:9] * 12) - 1:0] dccm_ext_in_pkt;
	input wire [(pt[909-:9] * 12) - 1:0] iccm_ext_in_pkt;
	input wire [pt[936-:9] - 1:1] iccm_rw_addr;
	input wire iccm_buf_correct_ecc;
	input wire iccm_correction_state;
	input wire iccm_wren;
	input wire iccm_rden;
	input wire [2:0] iccm_wr_size;
	input wire [77:0] iccm_wr_data;
	output wire [63:0] iccm_rd_data;
	output wire [77:0] iccm_rd_data_ecc;
	input wire [31:1] ic_rw_addr;
	input wire [pt[1060-:7] - 1:0] ic_tag_valid;
	input wire [pt[1060-:7] - 1:0] ic_wr_en;
	input wire ic_rd_en;
	input wire [63:0] ic_premux_data;
	input wire ic_sel_premux_data;
	input wire [((pt[1060-:7] * pt[1189-:7]) * 12) - 1:0] ic_data_ext_in_pkt;
	input wire [(pt[1060-:7] * 12) - 1:0] ic_tag_ext_in_pkt;
	input wire [(pt[1189-:7] * 71) - 1:0] ic_wr_data;
	input wire [70:0] ic_debug_wr_data;
	output wire [70:0] ic_debug_rd_data;
	input wire [pt[1104-:9]:3] ic_debug_addr;
	input wire ic_debug_rd_en;
	input wire ic_debug_wr_en;
	input wire ic_debug_tag_array;
	input wire [pt[1060-:7] - 1:0] ic_debug_way;
	output wire [63:0] ic_rd_data;
	output wire [25:0] ictag_debug_rd_data;
	output wire [pt[1189-:7] - 1:0] ic_eccerr;
	output wire [pt[1189-:7] - 1:0] ic_parerr;
	output wire [pt[1060-:7] - 1:0] ic_rd_hit;
	output wire ic_tag_perr;
	input wire scan_mode;
	wire active_clk;
	rvoclkhdr active_cg(
		.en(1'b1),
		.l1clk(active_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	generate
		if (pt[1365-:5] == 1) begin : Gen_dccm_enable
			eb1_lsu_dccm_mem #(.pt(pt)) dccm(
				.clk_override(dccm_clk_override),
				`ifdef USE_POWER_PINS
				.VPWR(VPWR),
				.VGND(VGND),
				`endif
				.clk(clk),
				.active_clk(active_clk),
				.rst_l(rst_l),
				.dccm_wren(dccm_wren),
				.dccm_rden(dccm_rden),
				.dccm_wr_addr_lo(dccm_wr_addr_lo),
				.dccm_wr_addr_hi(dccm_wr_addr_hi),
				.dccm_rd_addr_lo(dccm_rd_addr_lo),
				.dccm_rd_addr_hi(dccm_rd_addr_hi),
				.dccm_wr_data_lo(dccm_wr_data_lo),
				.dccm_wr_data_hi(dccm_wr_data_hi),
				.dccm_ext_in_pkt(dccm_ext_in_pkt),
				.dccm_rd_data_lo(dccm_rd_data_lo),
				.dccm_rd_data_hi(dccm_rd_data_hi),
				.scan_mode(scan_mode)
			);
		end
		else begin : Gen_dccm_disable
			assign dccm_rd_data_lo = {pt[1360-:10] {1'sb0}};
			assign dccm_rd_data_hi = {pt[1360-:10] {1'sb0}};
		end
	endgenerate
	generate
		if (pt[1120-:5]) begin : icache
			eb1_ifu_ic_mem #(.pt(pt)) icm(
				.clk_override(icm_clk_override),
				.*
			);
		end
		else begin
			assign ic_rd_hit[pt[1060-:7] - 1:0] = {pt[1060-:7] {1'sb0}};
			assign ic_tag_perr = 1'b0;
			assign ic_rd_data = {64 {1'sb0}};
			assign ictag_debug_rd_data = {26 {1'sb0}};
		end
	endgenerate
	generate
		if (pt[927-:5]) begin : iccm
			eb1_ifu_iccm_mem #(.pt(pt)) iccm(
				`ifdef USE_POWER_PINS
				.VPWR(VPWR),
				.VGND(VGND),
				`endif
				.clk(clk),
				.active_clk(active_clk),
				.rst_l(rst_l),
				.iccm_wren(iccm_wren),
				.iccm_rden(iccm_rden),
				.iccm_buf_correct_ecc(iccm_buf_correct_ecc),
				.iccm_correction_state(iccm_correction_state),
				.iccm_wr_size(iccm_wr_size),
				.iccm_wr_data(iccm_wr_data),
				.iccm_ext_in_pkt(iccm_ext_in_pkt),
				.iccm_rd_data_ecc(iccm_rd_data_ecc),
				.scan_mode(scan_mode),
				.clk_override(icm_clk_override),
				.iccm_rw_addr(iccm_rw_addr[pt[936-:9] - 1:1]),
				.iccm_rd_data(iccm_rd_data[63:0])
			);
		end
		else begin
			assign iccm_rd_data = {64 {1'sb0}};
			assign iccm_rd_data_ecc = {78 {1'sb0}};
		end
	endgenerate
endmodule
module eb1_pic_ctrl (
	clk,
	free_clk,
	rst_l,
	clk_override,
	io_clk_override,
	extintsrc_req,
	picm_rdaddr,
	picm_wraddr,
	picm_wr_data,
	picm_wren,
	picm_rden,
	picm_mken,
	meicurpl,
	meipt,
	mexintpend,
	claimid,
	pl,
	picm_rd_data,
	mhwakeup,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire free_clk;
	input wire rst_l;
	input wire clk_override;
	input wire io_clk_override;
	input wire [pt[44-:13] - 1:0] extintsrc_req;
	input wire [31:0] picm_rdaddr;
	input wire [31:0] picm_wraddr;
	input wire [31:0] picm_wr_data;
	input wire picm_wren;
	input wire picm_rden;
	input wire picm_mken;
	input wire [3:0] meicurpl;
	input wire [3:0] meipt;
	output wire mexintpend;
	output wire [7:0] claimid;
	output wire [3:0] pl;
	output wire [31:0] picm_rd_data;
	output wire mhwakeup;
	input wire scan_mode;
	localparam NUM_LEVELS = $clog2(pt[44-:13]);
	localparam INTPRIORITY_BASE_ADDR = pt[130-:36];
	localparam INTPEND_BASE_ADDR = pt[130-:36] + 32'h00001000;
	localparam INTENABLE_BASE_ADDR = pt[130-:36] + 32'h00002000;
	localparam EXT_INTR_PIC_CONFIG = pt[130-:36] + 32'h00003000;
	localparam EXT_INTR_GW_CONFIG = pt[130-:36] + 32'h00004000;
	localparam EXT_INTR_GW_CLEAR = pt[130-:36] + 32'h00005000;
	localparam INTPEND_SIZE = (pt[44-:13] < 32 ? 32 : (pt[44-:13] < 64 ? 64 : (pt[44-:13] < 128 ? 128 : (pt[44-:13] < 256 ? 256 : (pt[44-:13] < 512 ? 512 : 1024)))));
	localparam INT_GRPS = INTPEND_SIZE / 32;
	localparam INTPRIORITY_BITS = 4;
	localparam ID_BITS = 8;
	localparam signed [(pt[44-:13] * 32) - 1:0] GW_CONFIG = {pt[44-:13] {32'sd0}};
	localparam INT_ENABLE_GRPS = (pt[44-:13] - 1) / 4;
	wire [pt[44-:13] - 1:0] intenable_clk_enable;
	wire [INT_ENABLE_GRPS:0] intenable_clk_enable_grp;
	wire [INT_ENABLE_GRPS:0] gw_clk;
	wire addr_intpend_base_match;
	wire raddr_config_pic_match;
	wire raddr_intenable_base_match;
	wire raddr_intpriority_base_match;
	wire raddr_config_gw_base_match;
	wire waddr_config_pic_match;
	wire waddr_intpriority_base_match;
	wire waddr_intenable_base_match;
	wire waddr_config_gw_base_match;
	wire addr_clear_gw_base_match;
	wire mexintpend_in;
	wire mhwakeup_in;
	wire intpend_reg_read;
	wire [31:0] picm_rd_data_in;
	reg [31:0] intpend_rd_out;
	reg intenable_rd_out;
	reg [3:0] intpriority_rd_out;
	reg [1:0] gw_config_rd_out;
	wire [(pt[44-:13] * 4) - 1:0] intpriority_reg;
	wire [(pt[44-:13] * 4) - 1:0] intpriority_reg_inv;
	wire [pt[44-:13] - 1:0] intpriority_reg_we;
	wire [pt[44-:13] - 1:0] intpriority_reg_re;
	wire [(pt[44-:13] * 2) - 1:0] gw_config_reg;
	wire [pt[44-:13] - 1:0] intenable_reg;
	wire [pt[44-:13] - 1:0] intenable_reg_we;
	wire [pt[44-:13] - 1:0] intenable_reg_re;
	wire [pt[44-:13] - 1:0] gw_config_reg_we;
	wire [pt[44-:13] - 1:0] gw_config_reg_re;
	wire [pt[44-:13] - 1:0] gw_clear_reg_we;
	wire [INTPEND_SIZE - 1:0] intpend_reg_extended;
	wire [(pt[44-:13] * 4) - 1:0] intpend_w_prior_en;
	wire [(pt[44-:13] * 8) - 1:0] intpend_id;
	wire [3:0] maxint;
	wire [3:0] selected_int_priority;
	wire [(INT_GRPS * 32) - 1:0] intpend_rd_part_out;
	wire config_reg;
	wire intpriord;
	wire config_reg_we;
	wire config_reg_re;
	wire config_reg_in;
	wire prithresh_reg_write;
	wire prithresh_reg_read;
	wire intpriority_reg_read;
	wire intenable_reg_read;
	wire gw_config_reg_read;
	wire picm_wren_ff;
	wire picm_rden_ff;
	wire [31:0] picm_raddr_ff;
	wire [31:0] picm_waddr_ff;
	wire [31:0] picm_wr_data_ff;
	reg [3:0] mask;
	wire picm_mken_ff;
	wire [7:0] claimid_in;
	wire [3:0] pl_in;
	wire [3:0] pl_in_q;
	wire [pt[44-:13] - 1:0] extintsrc_req_sync;
	wire [pt[44-:13] - 1:0] extintsrc_req_gw;
	wire picm_bypass_ff;
	wire pic_raddr_c1_clken;
	wire pic_waddr_c1_clken;
	wire pic_data_c1_clken;
	wire pic_pri_c1_clken;
	wire pic_int_c1_clken;
	wire gw_config_c1_clken;
	wire pic_raddr_c1_clk;
	wire pic_data_c1_clk;
	wire pic_pri_c1_clk;
	wire pic_int_c1_clk;
	wire gw_config_c1_clk;
	assign pic_raddr_c1_clken = (picm_mken | picm_rden) | clk_override;
	assign pic_data_c1_clken = picm_wren | clk_override;
	assign pic_pri_c1_clken = ((waddr_intpriority_base_match & picm_wren_ff) | (raddr_intpriority_base_match & picm_rden_ff)) | clk_override;
	assign pic_int_c1_clken = ((waddr_intenable_base_match & picm_wren_ff) | (raddr_intenable_base_match & picm_rden_ff)) | clk_override;
	assign gw_config_c1_clken = ((waddr_config_gw_base_match & picm_wren_ff) | (raddr_config_gw_base_match & picm_rden_ff)) | clk_override;
	rvoclkhdr pic_addr_c1_cgc(
		.en(pic_raddr_c1_clken),
		.l1clk(pic_raddr_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr pic_data_c1_cgc(
		.en(pic_data_c1_clken),
		.l1clk(pic_data_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr pic_pri_c1_cgc(
		.en(pic_pri_c1_clken),
		.l1clk(pic_pri_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr pic_int_c1_cgc(
		.en(pic_int_c1_clken),
		.l1clk(pic_int_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr gw_config_c1_cgc(
		.en(gw_config_c1_clken),
		.l1clk(gw_config_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign raddr_intenable_base_match = picm_raddr_ff[31:NUM_LEVELS + 2] == INTENABLE_BASE_ADDR[31:NUM_LEVELS + 2];
	assign raddr_intpriority_base_match = picm_raddr_ff[31:NUM_LEVELS + 2] == INTPRIORITY_BASE_ADDR[31:NUM_LEVELS + 2];
	assign raddr_config_gw_base_match = picm_raddr_ff[31:NUM_LEVELS + 2] == EXT_INTR_GW_CONFIG[31:NUM_LEVELS + 2];
	assign raddr_config_pic_match = picm_raddr_ff[31:0] == EXT_INTR_PIC_CONFIG[31:0];
	assign addr_intpend_base_match = picm_raddr_ff[31:6] == INTPEND_BASE_ADDR[31:6];
	assign waddr_config_pic_match = picm_waddr_ff[31:0] == EXT_INTR_PIC_CONFIG[31:0];
	assign addr_clear_gw_base_match = picm_waddr_ff[31:NUM_LEVELS + 2] == EXT_INTR_GW_CLEAR[31:NUM_LEVELS + 2];
	assign waddr_intpriority_base_match = picm_waddr_ff[31:NUM_LEVELS + 2] == INTPRIORITY_BASE_ADDR[31:NUM_LEVELS + 2];
	assign waddr_intenable_base_match = picm_waddr_ff[31:NUM_LEVELS + 2] == INTENABLE_BASE_ADDR[31:NUM_LEVELS + 2];
	assign waddr_config_gw_base_match = picm_waddr_ff[31:NUM_LEVELS + 2] == EXT_INTR_GW_CONFIG[31:NUM_LEVELS + 2];
	assign picm_bypass_ff = (picm_rden_ff & picm_wren_ff) & (picm_raddr_ff[31:0] == picm_waddr_ff[31:0]);
	rvdff #(.WIDTH(32)) picm_radd_flop(
		.rst_l(rst_l),
		.din(picm_rdaddr),
		.dout(picm_raddr_ff),
		.clk(pic_raddr_c1_clk)
	);
	rvdff #(.WIDTH(32)) picm_wadd_flop(
		.rst_l(rst_l),
		.din(picm_wraddr),
		.dout(picm_waddr_ff),
		.clk(pic_data_c1_clk)
	);
	rvdff #(.WIDTH(1)) picm_wre_flop(
		.rst_l(rst_l),
		.din(picm_wren),
		.dout(picm_wren_ff),
		.clk(free_clk)
	);
	rvdff #(.WIDTH(1)) picm_rde_flop(
		.rst_l(rst_l),
		.din(picm_rden),
		.dout(picm_rden_ff),
		.clk(free_clk)
	);
	rvdff #(.WIDTH(1)) picm_mke_flop(
		.rst_l(rst_l),
		.din(picm_mken),
		.dout(picm_mken_ff),
		.clk(free_clk)
	);
	rvdff #(.WIDTH(32)) picm_dat_flop(
		.rst_l(rst_l),
		.din(picm_wr_data[31:0]),
		.dout(picm_wr_data_ff[31:0]),
		.clk(pic_data_c1_clk)
	);
	genvar p;
	generate
		for (p = 0; p <= INT_ENABLE_GRPS; p = p + 1) begin : IO_CLK_GRP
			if (p == INT_ENABLE_GRPS) begin : LAST_GRP
				assign intenable_clk_enable_grp[p] = |intenable_clk_enable[pt[44-:13] - 1:p * 4] | io_clk_override;
				rvoclkhdr intenable_c1_cgc(
					.en(intenable_clk_enable_grp[p]),
					.l1clk(gw_clk[p]),
					.clk(clk),
					.scan_mode(scan_mode)
				);
			end
			else begin : CLK_GRPS
				assign intenable_clk_enable_grp[p] = |intenable_clk_enable[(p * 4) + 3:p * 4] | io_clk_override;
				rvoclkhdr intenable_c1_cgc(
					.en(intenable_clk_enable_grp[p]),
					.l1clk(gw_clk[p]),
					.clk(clk),
					.scan_mode(scan_mode)
				);
			end
		end
	endgenerate
	genvar i;
	generate
		for (i = 0; i < pt[44-:13]; i = i + 1) begin : SETREG
			if (i > 0) begin : NON_ZERO_INT
				assign intpriority_reg_we[i] = (waddr_intpriority_base_match & (picm_waddr_ff[NUM_LEVELS + 1:2] == i)) & picm_wren_ff;
				assign intpriority_reg_re[i] = (raddr_intpriority_base_match & (picm_raddr_ff[NUM_LEVELS + 1:2] == i)) & picm_rden_ff;
				assign intenable_reg_we[i] = (waddr_intenable_base_match & (picm_waddr_ff[NUM_LEVELS + 1:2] == i)) & picm_wren_ff;
				assign intenable_reg_re[i] = (raddr_intenable_base_match & (picm_raddr_ff[NUM_LEVELS + 1:2] == i)) & picm_rden_ff;
				assign gw_config_reg_we[i] = (waddr_config_gw_base_match & (picm_waddr_ff[NUM_LEVELS + 1:2] == i)) & picm_wren_ff;
				assign gw_config_reg_re[i] = (raddr_config_gw_base_match & (picm_raddr_ff[NUM_LEVELS + 1:2] == i)) & picm_rden_ff;
				assign gw_clear_reg_we[i] = (addr_clear_gw_base_match & (picm_waddr_ff[NUM_LEVELS + 1:2] == i)) & picm_wren_ff;
				rvdffs #(.WIDTH(INTPRIORITY_BITS)) intpriority_ff(
					.rst_l(rst_l),
					.en(intpriority_reg_we[i]),
					.din(picm_wr_data_ff[3:0]),
					.dout(intpriority_reg[i * 4+:4]),
					.clk(pic_pri_c1_clk)
				);
				rvdffs #(.WIDTH(1)) intenable_ff(
					.rst_l(rst_l),
					.en(intenable_reg_we[i]),
					.din(picm_wr_data_ff[0]),
					.dout(intenable_reg[i]),
					.clk(pic_int_c1_clk)
				);
				assign intenable_clk_enable[i] = ((gw_config_reg[(i * 2) + 1] | intenable_reg_we[i]) | intenable_reg[i]) | gw_clear_reg_we[i];
				rvsyncss_fpga #(.WIDTH(1)) sync_inst(
					.gw_clk(gw_clk[i / 4]),
					.rawclk(clk),
					.clken(intenable_clk_enable_grp[i / 4]),
					.dout(extintsrc_req_sync[i]),
					.din(extintsrc_req[i]),
					.rst_l(rst_l)
				);
				rvdffs #(.WIDTH(2)) gw_config_ff(
					.rst_l(rst_l),
					.en(gw_config_reg_we[i]),
					.din(picm_wr_data_ff[1:0]),
					.dout(gw_config_reg[i * 2+:2]),
					.clk(gw_config_c1_clk)
				);
				eb1_configurable_gw config_gw_inst(
					.rst_l(rst_l),
					.gw_clk(gw_clk[i / 4]),
					.rawclk(clk),
					.clken(intenable_clk_enable_grp[i / 4]),
					.extintsrc_req_sync(extintsrc_req_sync[i]),
					.meigwctrl_polarity(gw_config_reg[i * 2]),
					.meigwctrl_type(gw_config_reg[(i * 2) + 1]),
					.meigwclr(gw_clear_reg_we[i]),
					.extintsrc_req_config(extintsrc_req_gw[i])
				);
			end
			else begin : INT_ZERO
				assign intpriority_reg_we[i] = 1'b0;
				assign intpriority_reg_re[i] = 1'b0;
				assign intenable_reg_we[i] = 1'b0;
				assign intenable_reg_re[i] = 1'b0;
				assign gw_config_reg_we[i] = 1'b0;
				assign gw_config_reg_re[i] = 1'b0;
				assign gw_clear_reg_we[i] = 1'b0;
				assign gw_config_reg[i * 2+:2] = {2 {1'sb0}};
				assign intpriority_reg[i * 4+:4] = {INTPRIORITY_BITS {1'b0}};
				assign intenable_reg[i] = 1'b0;
				assign extintsrc_req_gw[i] = 1'b0;
				assign extintsrc_req_sync[i] = 1'b0;
				assign intenable_clk_enable[i] = 1'b0;
			end
			assign intpriority_reg_inv[i * 4+:4] = (intpriord ? ~intpriority_reg[i * 4+:4] : intpriority_reg[i * 4+:4]);
			assign intpend_w_prior_en[i * 4+:4] = {INTPRIORITY_BITS {extintsrc_req_gw[i] & intenable_reg[i]}} & intpriority_reg_inv[i * 4+:4];
			assign intpend_id[i * 8+:8] = i;
		end
	endgenerate
	assign pl_in[3:0] = selected_int_priority[3:0];
	genvar l;
	genvar m;
	genvar j;
	genvar k;
	generate
		if (pt[135-:5] == 1) begin : genblock
			wire [(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))))) + 1) * 4) + ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) * 4) - 1) : (((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1)))) + 1) * 4) + ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) * 4) - 1)):(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) * 4 : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) * 4)] level_intpend_w_prior_en;
			wire [(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))))) + 1) * 8) + ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) * 8) - 1) : (((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1)))) + 1) * 8) + ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) * 8) - 1)):(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) * 8 : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) * 8)] level_intpend_id;
			wire [((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))))) + 1) * 4) + (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) * 4) - 1) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)))) + 1) * 4) + (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) * 4) - 1)):((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) * 4 : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) * 4)] levelx_intpend_w_prior_en;
			wire [((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))))) + 1) * 8) + (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) * 8) - 1) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)))) + 1) * 8) + (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) * 8) - 1)):((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) * 8 : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) * 8)] levelx_intpend_id;
			assign level_intpend_w_prior_en[4 * (((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) - (((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2)) - 1) : ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) - (((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2)) - 1) : ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1)))))+:4 * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))] = {12'b000000000000, intpend_w_prior_en[4 * ((pt[44-:13] - 1) - (pt[44-:13] - 1))+:4 * pt[44-:13]]};
			assign level_intpend_id[8 * (((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) - (((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2)) - 1) : ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - ((((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) - (((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2)) - 1) : ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) : (((((NUM_LEVELS / 2) >= 0 ? 0 : NUM_LEVELS / 2) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1) : (pt[44-:13] + 2) - ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 2 : ((pt[44-:13] + 2) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1))) + ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) - 1)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1)))))+:8 * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))] = {24'b000000000000000000000000, intpend_id[8 * ((pt[44-:13] - 1) - (pt[44-:13] - 1))+:8 * pt[44-:13]]};
			wire [((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) * 4) - 1 : ((1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) * 4) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) * 4) - 1)):((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) * 4)] l2_intpend_w_prior_en_ff;
			wire [((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) * 8) - 1 : ((1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) * 8) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) * 8) - 1)):((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) * 8)] l2_intpend_id_ff;
			assign levelx_intpend_w_prior_en[4 * ((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) - ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - 1) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) - ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - 1) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)))))+:4 * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))] = {{4 {1'b0}}, l2_intpend_w_prior_en_ff[4 * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1)) : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1)))+:4 * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))]};
			assign levelx_intpend_id[8 * ((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) - ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - 1) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - (((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) - ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - 1) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) : ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - ((NUM_LEVELS / 2) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) - 1)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)))))+:8 * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))] = {{8 {1'b1}}, l2_intpend_id_ff[8 * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1)) : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1) - (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2)))) - 1) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? pt[44-:13] / (2 ** (NUM_LEVELS / 2)) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))) - 1)))+:8 * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1 : 1 - (pt[44-:13] / (2 ** (NUM_LEVELS / 2))))]};
			for (l = 0; l < (NUM_LEVELS / 2); l = l + 1) begin : TOP_LEVEL
				for (m = 0; m <= (pt[44-:13] / (2 ** (l + 1))); m = m + 1) begin : COMPARE
					if (m == (pt[44-:13] / (2 ** (l + 1)))) begin
						assign level_intpend_w_prior_en[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m + 1 : (pt[44-:13] + 2) - (m + 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m + 1 : (pt[44-:13] + 2) - (m + 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 4+:4] = {4 {1'sb0}};
						assign level_intpend_id[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m + 1 : (pt[44-:13] + 2) - (m + 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m + 1 : (pt[44-:13] + 2) - (m + 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 8+:8] = {8 {1'sb0}};
					end
					eb1_cmp_and_mux #(
						.ID_BITS(ID_BITS),
						.INTPRIORITY_BITS(INTPRIORITY_BITS)
					) cmp_l1(
						.a_id(level_intpend_id[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? 2 * m : (pt[44-:13] + 2) - (2 * m)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? 2 * m : (pt[44-:13] + 2) - (2 * m))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 8+:8]),
						.a_priority(level_intpend_w_prior_en[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? 2 * m : (pt[44-:13] + 2) - (2 * m)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? 2 * m : (pt[44-:13] + 2) - (2 * m))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 4+:4]),
						.b_id(level_intpend_id[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 2) - ((2 * m) + 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 2) - ((2 * m) + 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 8+:8]),
						.b_priority(level_intpend_w_prior_en[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 2) - ((2 * m) + 1)) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l : (NUM_LEVELS / 2) - l) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 2) - ((2 * m) + 1))) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 4+:4]),
						.out_id(level_intpend_id[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m : (pt[44-:13] + 2) - m) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m : (pt[44-:13] + 2) - m)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 8+:8]),
						.out_priority(level_intpend_w_prior_en[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m : (pt[44-:13] + 2) - m) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? l + 1 : (NUM_LEVELS / 2) - (l + 1)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? m : (pt[44-:13] + 2) - m)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 4+:4])
					);
				end
			end
			for (i = 0; i <= (pt[44-:13] / (2 ** (NUM_LEVELS / 2))); i = i + 1) begin : MIDDLE_FLOPS
				rvdff #(.WIDTH(INTPRIORITY_BITS)) leveb1_intpend_prior_reg(
					.rst_l(rst_l),
					.din(level_intpend_w_prior_en[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - (NUM_LEVELS / 2)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? i : (pt[44-:13] + 2) - i) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - (NUM_LEVELS / 2)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? i : (pt[44-:13] + 2) - i)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 4+:4]),
					.dout(l2_intpend_w_prior_en_ff[((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? i : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) - i) * 4+:4]),
					.clk(free_clk)
				);
				rvdff #(.WIDTH(ID_BITS)) leveb1_intpend_id_reg(
					.rst_l(rst_l),
					.din(level_intpend_id[(((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))) >= ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) ? (((NUM_LEVELS / 2) >= 0 ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - (NUM_LEVELS / 2)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? i : (pt[44-:13] + 2) - i) : ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? 0 : pt[44-:13] + 2) : ((pt[44-:13] + 2) >= 0 ? (NUM_LEVELS / 2) * (pt[44-:13] + 3) : (pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2))))) - (((((NUM_LEVELS / 2) >= 0 ? NUM_LEVELS / 2 : (NUM_LEVELS / 2) - (NUM_LEVELS / 2)) * ((pt[44-:13] + 2) >= 0 ? pt[44-:13] + 3 : 1 - (pt[44-:13] + 2))) + ((pt[44-:13] + 2) >= 0 ? i : (pt[44-:13] + 2) - i)) - ((NUM_LEVELS / 2) >= 0 ? ((pt[44-:13] + 2) >= 0 ? (((NUM_LEVELS / 2) + 1) * (pt[44-:13] + 3)) - 1 : (((NUM_LEVELS / 2) + 1) * (1 - (pt[44-:13] + 2))) + (pt[44-:13] + 1)) : ((pt[44-:13] + 2) >= 0 ? ((1 - (NUM_LEVELS / 2)) * (pt[44-:13] + 3)) + (((NUM_LEVELS / 2) * (pt[44-:13] + 3)) - 1) : ((1 - (NUM_LEVELS / 2)) * (1 - (pt[44-:13] + 2))) + (((pt[44-:13] + 2) + ((NUM_LEVELS / 2) * (1 - (pt[44-:13] + 2)))) - 1))))) * 8+:8]),
					.dout(l2_intpend_id_ff[((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) >= 0 ? i : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) - i) * 8+:8]),
					.clk(free_clk)
				);
			end
			for (j = NUM_LEVELS / 2; j < NUM_LEVELS; j = j + 1) begin : BOT_LEVELS
				for (k = 0; k <= (pt[44-:13] / (2 ** (j + 1))); k = k + 1) begin : COMPARE
					if (k == (pt[44-:13] / (2 ** (j + 1)))) begin
						assign levelx_intpend_w_prior_en[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (k + 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (k + 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 4+:4] = {4 {1'sb0}};
						assign levelx_intpend_id[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (k + 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (k + 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 8+:8] = {8 {1'sb0}};
					end
					eb1_cmp_and_mux #(
						.ID_BITS(ID_BITS),
						.INTPRIORITY_BITS(INTPRIORITY_BITS)
					) cmp_l1(
						.a_id(levelx_intpend_id[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 2 * k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (2 * k)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 2 * k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (2 * k))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 8+:8]),
						.a_priority(levelx_intpend_w_prior_en[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 2 * k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (2 * k)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 2 * k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - (2 * k))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 4+:4]),
						.b_id(levelx_intpend_id[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (2 * k) + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - ((2 * k) + 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (2 * k) + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - ((2 * k) + 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 8+:8]),
						.b_priority(levelx_intpend_w_prior_en[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (2 * k) + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - ((2 * k) + 1)) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j : (NUM_LEVELS / 2) - (j - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (2 * k) + 1 : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - ((2 * k) + 1))) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 4+:4]),
						.out_id(levelx_intpend_id[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - k) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - k)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 8+:8]),
						.out_priority(levelx_intpend_w_prior_en[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - k) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? j + 1 : (NUM_LEVELS / 2) - ((j + 1) - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? k : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) - k)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 4+:4])
					);
				end
			end
			assign claimid_in[7:0] = levelx_intpend_id[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS : (NUM_LEVELS / 2) - (NUM_LEVELS - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS : (NUM_LEVELS / 2) - (NUM_LEVELS - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 8+:8];
			assign selected_int_priority[3:0] = levelx_intpend_w_prior_en[((NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))) >= (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) ? ((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS : (NUM_LEVELS / 2) - (NUM_LEVELS - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) : (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2) : ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))))) - ((((NUM_LEVELS >= (NUM_LEVELS / 2) ? NUM_LEVELS : (NUM_LEVELS / 2) - (NUM_LEVELS - NUM_LEVELS)) * (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2 : 1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? 0 : (pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)) - (NUM_LEVELS >= (NUM_LEVELS / 2) ? (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + (((NUM_LEVELS / 2) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : (((NUM_LEVELS - (NUM_LEVELS / 2)) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + ((NUM_LEVELS / 2) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1)) : (((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) >= 0 ? ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) + ((NUM_LEVELS * ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 2)) - 1) : ((((NUM_LEVELS / 2) - NUM_LEVELS) + 1) * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1))) + ((((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1) + (NUM_LEVELS * (1 - ((pt[44-:13] / (2 ** (NUM_LEVELS / 2))) + 1)))) - 1))))) * 4+:4];
		end
		else begin : genblock
			wire [((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))))) + 1) * 4) + (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) * 4) - 1) : ((((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1)))) + 1) * 4) + (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) * 4) - 1)):((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) * 4 : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) * 4)] level_intpend_w_prior_en;
			wire [((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))))) + 1) * 8) + (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) * 8) - 1) : ((((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1)))) + 1) * 8) + (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) * 8) - 1)):((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) * 8 : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) * 8)] level_intpend_id;
			assign level_intpend_w_prior_en[4 * ((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) - (((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1)) - 1) : ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) - (((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1)) - 1) : ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1)))))+:4 * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))] = {{8 {1'b0}}, intpend_w_prior_en[4 * ((pt[44-:13] - 1) - (pt[44-:13] - 1))+:4 * pt[44-:13]]};
			assign level_intpend_id[8 * ((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) - (((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1)) - 1) : ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - (((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) - (((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1)) - 1) : ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) : ((((NUM_LEVELS >= 0 ? 0 : NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1) : (pt[44-:13] + 1) - ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 1 : ((pt[44-:13] + 1) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1))) + ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) - 1)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1)))))+:8 * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))] = {{16 {1'b1}}, intpend_id[8 * ((pt[44-:13] - 1) - (pt[44-:13] - 1))+:8 * pt[44-:13]]};
			for (l = 0; l < NUM_LEVELS; l = l + 1) begin : LEVEL
				for (m = 0; m <= (pt[44-:13] / (2 ** (l + 1))); m = m + 1) begin : COMPARE
					if (m == (pt[44-:13] / (2 ** (l + 1)))) begin
						assign level_intpend_w_prior_en[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m + 1 : (pt[44-:13] + 1) - (m + 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m + 1 : (pt[44-:13] + 1) - (m + 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 4+:4] = {4 {1'sb0}};
						assign level_intpend_id[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m + 1 : (pt[44-:13] + 1) - (m + 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m + 1 : (pt[44-:13] + 1) - (m + 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 8+:8] = {8 {1'sb0}};
					end
					eb1_cmp_and_mux #(
						.ID_BITS(ID_BITS),
						.INTPRIORITY_BITS(INTPRIORITY_BITS)
					) cmp_l1(
						.a_id(level_intpend_id[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 2 * m : (pt[44-:13] + 1) - (2 * m)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 2 * m : (pt[44-:13] + 1) - (2 * m))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 8+:8]),
						.a_priority(level_intpend_w_prior_en[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 2 * m : (pt[44-:13] + 1) - (2 * m)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 2 * m : (pt[44-:13] + 1) - (2 * m))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 4+:4]),
						.b_id(level_intpend_id[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 1) - ((2 * m) + 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 1) - ((2 * m) + 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 8+:8]),
						.b_priority(level_intpend_w_prior_en[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 1) - ((2 * m) + 1)) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l : NUM_LEVELS - l) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? (2 * m) + 1 : (pt[44-:13] + 1) - ((2 * m) + 1))) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 4+:4]),
						.out_id(level_intpend_id[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m : (pt[44-:13] + 1) - m) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m : (pt[44-:13] + 1) - m)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 8+:8]),
						.out_priority(level_intpend_w_prior_en[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m : (pt[44-:13] + 1) - m) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? l + 1 : NUM_LEVELS - (l + 1)) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? m : (pt[44-:13] + 1) - m)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 4+:4])
					);
				end
			end
			assign claimid_in[7:0] = level_intpend_id[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? NUM_LEVELS : NUM_LEVELS - NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? NUM_LEVELS : NUM_LEVELS - NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 8+:8];
			assign selected_int_priority[3:0] = level_intpend_w_prior_en[((NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))) >= (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) ? ((NUM_LEVELS >= 0 ? NUM_LEVELS : NUM_LEVELS - NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1) : ((pt[44-:13] + 1) >= 0 ? NUM_LEVELS * (pt[44-:13] + 2) : (pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1))))) - ((((NUM_LEVELS >= 0 ? NUM_LEVELS : NUM_LEVELS - NUM_LEVELS) * ((pt[44-:13] + 1) >= 0 ? pt[44-:13] + 2 : 1 - (pt[44-:13] + 1))) + ((pt[44-:13] + 1) >= 0 ? 0 : pt[44-:13] + 1)) - (NUM_LEVELS >= 0 ? ((pt[44-:13] + 1) >= 0 ? ((NUM_LEVELS + 1) * (pt[44-:13] + 2)) - 1 : ((NUM_LEVELS + 1) * (1 - (pt[44-:13] + 1))) + pt[44-:13]) : ((pt[44-:13] + 1) >= 0 ? ((1 - NUM_LEVELS) * (pt[44-:13] + 2)) + ((NUM_LEVELS * (pt[44-:13] + 2)) - 1) : ((1 - NUM_LEVELS) * (1 - (pt[44-:13] + 1))) + (((pt[44-:13] + 1) + (NUM_LEVELS * (1 - (pt[44-:13] + 1)))) - 1))))) * 4+:4];
		end
	endgenerate
	assign config_reg_we = waddr_config_pic_match & picm_wren_ff;
	assign config_reg_re = raddr_config_pic_match & picm_rden_ff;
	assign config_reg_in = picm_wr_data_ff[0];
	rvdffs #(.WIDTH(1)) config_reg_ff(
		.rst_l(rst_l),
		.clk(free_clk),
		.en(config_reg_we),
		.din(config_reg_in),
		.dout(config_reg)
	);
	assign intpriord = config_reg;
	assign pl_in_q[3:0] = (intpriord ? ~pl_in : pl_in);
	rvdff #(.WIDTH(ID_BITS)) claimid_ff(
		.rst_l(rst_l),
		.din(claimid_in[7:0]),
		.dout(claimid[7:0]),
		.clk(free_clk)
	);
	rvdff #(.WIDTH(INTPRIORITY_BITS)) pl_ff(
		.rst_l(rst_l),
		.din(pl_in_q[3:0]),
		.dout(pl[3:0]),
		.clk(free_clk)
	);
	wire [3:0] meipt_inv;
	wire [3:0] meicurpl_inv;
	assign meipt_inv[3:0] = (intpriord ? ~meipt[3:0] : meipt[3:0]);
	assign meicurpl_inv[3:0] = (intpriord ? ~meicurpl[3:0] : meicurpl[3:0]);
	assign mexintpend_in = (selected_int_priority[3:0] > meipt_inv[3:0]) & (selected_int_priority[3:0] > meicurpl_inv[3:0]);
	rvdff #(.WIDTH(1)) mexintpend_ff(
		.rst_l(rst_l),
		.clk(free_clk),
		.din(mexintpend_in),
		.dout(mexintpend)
	);
	assign maxint[3:0] = (intpriord ? 0 : 15);
	assign mhwakeup_in = pl_in_q[3:0] == maxint;
	rvdff #(.WIDTH(1)) wake_up_ff(
		.rst_l(rst_l),
		.clk(free_clk),
		.din(mhwakeup_in),
		.dout(mhwakeup)
	);
	assign intpend_reg_read = addr_intpend_base_match & picm_rden_ff;
	assign intpriority_reg_read = raddr_intpriority_base_match & picm_rden_ff;
	assign intenable_reg_read = raddr_intenable_base_match & picm_rden_ff;
	assign gw_config_reg_read = raddr_config_gw_base_match & picm_rden_ff;
	assign intpend_reg_extended[INTPEND_SIZE - 1:0] = {{INTPEND_SIZE - pt[44-:13] {1'b0}}, extintsrc_req_gw[pt[44-:13] - 1:0]};
	generate
		for (i = 0; i < INT_GRPS; i = i + 1) assign intpend_rd_part_out[i * 32+:32] = {32 {intpend_reg_read & (picm_raddr_ff[5:2] == i)}} & intpend_reg_extended[(32 * i) + 31:32 * i];
	endgenerate
	always @(*) begin : INTPEND_RD
		intpend_rd_out = {32 {1'sb0}};
		begin : sv2v_autoblock_34
			reg signed [31:0] i;
			for (i = 0; i < INT_GRPS; i = i + 1)
				intpend_rd_out = intpend_rd_out | intpend_rd_part_out[i * 32+:32];
		end
	end
	always @(*) begin : INTEN_RD
		intenable_rd_out = 1'b0;
		intpriority_rd_out = {4 {1'sb0}};
		gw_config_rd_out = {2 {1'sb0}};
		begin : sv2v_autoblock_35
			reg signed [31:0] i;
			for (i = 0; i < pt[44-:13]; i = i + 1)
				begin
					if (intenable_reg_re[i])
						intenable_rd_out = intenable_reg[i];
					if (intpriority_reg_re[i])
						intpriority_rd_out = intpriority_reg[i * 4+:4];
					if (gw_config_reg_re[i])
						gw_config_rd_out = gw_config_reg[i * 2+:2];
				end
		end
	end
	assign picm_rd_data_in[31:0] = (((((((({32 {intpend_reg_read}} & intpend_rd_out) | ({32 {intpriority_reg_read}} & {{28 {1'b0}}, intpriority_rd_out})) | ({32 {intenable_reg_read}} & {31'b0000000000000000000000000000000, intenable_rd_out})) | ({32 {gw_config_reg_read}} & {30'b000000000000000000000000000000, gw_config_rd_out})) | ({32 {config_reg_re}} & {31'b0000000000000000000000000000000, config_reg})) | ({32 {picm_mken_ff & mask[3]}} & 32'b00000000000000000000000000000011)) | ({32 {picm_mken_ff & mask[2]}} & 32'b00000000000000000000000000000001)) | ({32 {picm_mken_ff & mask[1]}} & 32'b00000000000000000000000000001111)) | ({32 {picm_mken_ff & mask[0]}} & 32'b00000000000000000000000000000000);
	assign picm_rd_data[31:0] = (picm_bypass_ff ? picm_wr_data_ff[31:0] : picm_rd_data_in[31:0]);
	wire [14:0] address;
	assign address[14:0] = picm_raddr_ff[14:0];
	always @(*)
		case (address[14:0])
			15'b011000000000000: mask[3:0] = 4'b0100;
			15'b100000000000100: mask[3:0] = 4'b1000;
			15'b100000000001000: mask[3:0] = 4'b1000;
			15'b100000000001100: mask[3:0] = 4'b1000;
			15'b100000000010000: mask[3:0] = 4'b1000;
			15'b100000000010100: mask[3:0] = 4'b1000;
			15'b100000000011000: mask[3:0] = 4'b1000;
			15'b100000000011100: mask[3:0] = 4'b1000;
			15'b100000000100000: mask[3:0] = 4'b1000;
			15'b100000000100100: mask[3:0] = 4'b1000;
			15'b100000000101000: mask[3:0] = 4'b1000;
			15'b100000000101100: mask[3:0] = 4'b1000;
			15'b100000000110000: mask[3:0] = 4'b1000;
			15'b100000000110100: mask[3:0] = 4'b1000;
			15'b100000000111000: mask[3:0] = 4'b1000;
			15'b100000000111100: mask[3:0] = 4'b1000;
			15'b100000001000000: mask[3:0] = 4'b1000;
			15'b100000001000100: mask[3:0] = 4'b1000;
			15'b100000001001000: mask[3:0] = 4'b1000;
			15'b100000001001100: mask[3:0] = 4'b1000;
			15'b100000001010000: mask[3:0] = 4'b1000;
			15'b100000001010100: mask[3:0] = 4'b1000;
			15'b100000001011000: mask[3:0] = 4'b1000;
			15'b100000001011100: mask[3:0] = 4'b1000;
			15'b100000001100000: mask[3:0] = 4'b1000;
			15'b100000001100100: mask[3:0] = 4'b1000;
			15'b100000001101000: mask[3:0] = 4'b1000;
			15'b100000001101100: mask[3:0] = 4'b1000;
			15'b100000001110000: mask[3:0] = 4'b1000;
			15'b100000001110100: mask[3:0] = 4'b1000;
			15'b100000001111000: mask[3:0] = 4'b1000;
			15'b100000001111100: mask[3:0] = 4'b1000;
			15'b010000000000100: mask[3:0] = 4'b0100;
			15'b010000000001000: mask[3:0] = 4'b0100;
			15'b010000000001100: mask[3:0] = 4'b0100;
			15'b010000000010000: mask[3:0] = 4'b0100;
			15'b010000000010100: mask[3:0] = 4'b0100;
			15'b010000000011000: mask[3:0] = 4'b0100;
			15'b010000000011100: mask[3:0] = 4'b0100;
			15'b010000000100000: mask[3:0] = 4'b0100;
			15'b010000000100100: mask[3:0] = 4'b0100;
			15'b010000000101000: mask[3:0] = 4'b0100;
			15'b010000000101100: mask[3:0] = 4'b0100;
			15'b010000000110000: mask[3:0] = 4'b0100;
			15'b010000000110100: mask[3:0] = 4'b0100;
			15'b010000000111000: mask[3:0] = 4'b0100;
			15'b010000000111100: mask[3:0] = 4'b0100;
			15'b010000001000000: mask[3:0] = 4'b0100;
			15'b010000001000100: mask[3:0] = 4'b0100;
			15'b010000001001000: mask[3:0] = 4'b0100;
			15'b010000001001100: mask[3:0] = 4'b0100;
			15'b010000001010000: mask[3:0] = 4'b0100;
			15'b010000001010100: mask[3:0] = 4'b0100;
			15'b010000001011000: mask[3:0] = 4'b0100;
			15'b010000001011100: mask[3:0] = 4'b0100;
			15'b010000001100000: mask[3:0] = 4'b0100;
			15'b010000001100100: mask[3:0] = 4'b0100;
			15'b010000001101000: mask[3:0] = 4'b0100;
			15'b010000001101100: mask[3:0] = 4'b0100;
			15'b010000001110000: mask[3:0] = 4'b0100;
			15'b010000001110100: mask[3:0] = 4'b0100;
			15'b010000001111000: mask[3:0] = 4'b0100;
			15'b010000001111100: mask[3:0] = 4'b0100;
			15'b000000000000100: mask[3:0] = 4'b0010;
			15'b000000000001000: mask[3:0] = 4'b0010;
			15'b000000000001100: mask[3:0] = 4'b0010;
			15'b000000000010000: mask[3:0] = 4'b0010;
			15'b000000000010100: mask[3:0] = 4'b0010;
			15'b000000000011000: mask[3:0] = 4'b0010;
			15'b000000000011100: mask[3:0] = 4'b0010;
			15'b000000000100000: mask[3:0] = 4'b0010;
			15'b000000000100100: mask[3:0] = 4'b0010;
			15'b000000000101000: mask[3:0] = 4'b0010;
			15'b000000000101100: mask[3:0] = 4'b0010;
			15'b000000000110000: mask[3:0] = 4'b0010;
			15'b000000000110100: mask[3:0] = 4'b0010;
			15'b000000000111000: mask[3:0] = 4'b0010;
			15'b000000000111100: mask[3:0] = 4'b0010;
			15'b000000001000000: mask[3:0] = 4'b0010;
			15'b000000001000100: mask[3:0] = 4'b0010;
			15'b000000001001000: mask[3:0] = 4'b0010;
			15'b000000001001100: mask[3:0] = 4'b0010;
			15'b000000001010000: mask[3:0] = 4'b0010;
			15'b000000001010100: mask[3:0] = 4'b0010;
			15'b000000001011000: mask[3:0] = 4'b0010;
			15'b000000001011100: mask[3:0] = 4'b0010;
			15'b000000001100000: mask[3:0] = 4'b0010;
			15'b000000001100100: mask[3:0] = 4'b0010;
			15'b000000001101000: mask[3:0] = 4'b0010;
			15'b000000001101100: mask[3:0] = 4'b0010;
			15'b000000001110000: mask[3:0] = 4'b0010;
			15'b000000001110100: mask[3:0] = 4'b0010;
			15'b000000001111000: mask[3:0] = 4'b0010;
			15'b000000001111100: mask[3:0] = 4'b0010;
			default: mask[3:0] = 4'b0001;
		endcase
endmodule
module eb1_cmp_and_mux (
	a_id,
	a_priority,
	b_id,
	b_priority,
	out_id,
	out_priority
);
	parameter ID_BITS = 8;
	parameter INTPRIORITY_BITS = 4;
	input wire [ID_BITS - 1:0] a_id;
	input wire [INTPRIORITY_BITS - 1:0] a_priority;
	input wire [ID_BITS - 1:0] b_id;
	input wire [INTPRIORITY_BITS - 1:0] b_priority;
	output wire [ID_BITS - 1:0] out_id;
	output wire [INTPRIORITY_BITS - 1:0] out_priority;
	wire a_is_lt_b;
	assign a_is_lt_b = a_priority[INTPRIORITY_BITS - 1:0] < b_priority[INTPRIORITY_BITS - 1:0];
	assign out_id[ID_BITS - 1:0] = (a_is_lt_b ? b_id[ID_BITS - 1:0] : a_id[ID_BITS - 1:0]);
	assign out_priority[INTPRIORITY_BITS - 1:0] = (a_is_lt_b ? b_priority[INTPRIORITY_BITS - 1:0] : a_priority[INTPRIORITY_BITS - 1:0]);
endmodule
module eb1_configurable_gw (
	gw_clk,
	rawclk,
	clken,
	rst_l,
	extintsrc_req_sync,
	meigwctrl_polarity,
	meigwctrl_type,
	meigwclr,
	extintsrc_req_config
);
	input wire gw_clk;
	input wire rawclk;
	input wire clken;
	input wire rst_l;
	input wire extintsrc_req_sync;
	input wire meigwctrl_polarity;
	input wire meigwctrl_type;
	input wire meigwclr;
	output wire extintsrc_req_config;
	wire gw_int_pending_in;
	wire gw_int_pending;
	assign gw_int_pending_in = (extintsrc_req_sync ^ meigwctrl_polarity) | (gw_int_pending & ~meigwclr);
	rvdff_fpga #(.WIDTH(1)) int_pend_ff(
		.rst_l(rst_l),
		.clk(gw_clk),
		.rawclk(rawclk),
		.clken(clken),
		.din(gw_int_pending_in),
		.dout(gw_int_pending)
	);
	assign extintsrc_req_config = (meigwctrl_type ? (extintsrc_req_sync ^ meigwctrl_polarity) | gw_int_pending : extintsrc_req_sync ^ meigwctrl_polarity);
endmodule
module ahb_to_axi4 (
	clk,
	rst_l,
	scan_mode,
	bus_clk_en,
	clk_override,
	axi_awvalid,
	axi_awready,
	axi_awid,
	axi_awaddr,
	axi_awsize,
	axi_awprot,
	axi_awlen,
	axi_awburst,
	axi_wvalid,
	axi_wready,
	axi_wdata,
	axi_wstrb,
	axi_wlast,
	axi_bvalid,
	axi_bready,
	axi_bresp,
	axi_bid,
	axi_arvalid,
	axi_arready,
	axi_arid,
	axi_araddr,
	axi_arsize,
	axi_arprot,
	axi_arlen,
	axi_arburst,
	axi_rvalid,
	axi_rready,
	axi_rid,
	axi_rdata,
	axi_rresp,
	ahb_haddr,
	ahb_hburst,
	ahb_hmastlock,
	ahb_hprot,
	ahb_hsize,
	ahb_htrans,
	ahb_hwrite,
	ahb_hwdata,
	ahb_hsel,
	ahb_hreadyin,
	ahb_hrdata,
	ahb_hreadyout,
	ahb_hresp
);
	parameter TAG = 1;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input clk;
	input rst_l;
	input scan_mode;
	input bus_clk_en;
	input clk_override;
	output wire axi_awvalid;
	input wire axi_awready;
	output wire [TAG - 1:0] axi_awid;
	output wire [31:0] axi_awaddr;
	output wire [2:0] axi_awsize;
	output wire [2:0] axi_awprot;
	output wire [7:0] axi_awlen;
	output wire [1:0] axi_awburst;
	output wire axi_wvalid;
	input wire axi_wready;
	output wire [63:0] axi_wdata;
	output wire [7:0] axi_wstrb;
	output wire axi_wlast;
	input wire axi_bvalid;
	output wire axi_bready;
	input wire [1:0] axi_bresp;
	input wire [TAG - 1:0] axi_bid;
	output wire axi_arvalid;
	input wire axi_arready;
	output wire [TAG - 1:0] axi_arid;
	output wire [31:0] axi_araddr;
	output wire [2:0] axi_arsize;
	output wire [2:0] axi_arprot;
	output wire [7:0] axi_arlen;
	output wire [1:0] axi_arburst;
	input wire axi_rvalid;
	output wire axi_rready;
	input wire [TAG - 1:0] axi_rid;
	input wire [63:0] axi_rdata;
	input wire [1:0] axi_rresp;
	input wire [31:0] ahb_haddr;
	input wire [2:0] ahb_hburst;
	input wire ahb_hmastlock;
	input wire [3:0] ahb_hprot;
	input wire [2:0] ahb_hsize;
	input wire [1:0] ahb_htrans;
	input wire ahb_hwrite;
	input wire [63:0] ahb_hwdata;
	input wire ahb_hsel;
	input wire ahb_hreadyin;
	output wire [63:0] ahb_hrdata;
	output wire ahb_hreadyout;
	output wire ahb_hresp;
	wire [7:0] master_wstrb;
	wire [1:0] buf_state;
	reg [1:0] buf_nxtstate;
	reg buf_state_en;
	reg buf_read_error_in;
	wire buf_read_error;
	wire [63:0] buf_rdata;
	wire ahb_hready;
	wire ahb_hready_q;
	wire [1:0] ahb_htrans_in;
	wire [1:0] ahb_htrans_q;
	wire [2:0] ahb_hsize_q;
	wire ahb_hwrite_q;
	wire [31:0] ahb_haddr_q;
	wire [63:0] ahb_hwdata_q;
	wire ahb_hresp_q;
	wire ahb_addr_in_dccm;
	wire ahb_addr_in_iccm;
	wire ahb_addr_in_pic;
	wire ahb_addr_in_dccm_region_nc;
	wire ahb_addr_in_iccm_region_nc;
	wire ahb_addr_in_pic_region_nc;
	reg buf_rdata_en;
	wire ahb_addr_clk_en;
	wire buf_rdata_clk_en;
	wire bus_clk;
	wire ahb_addr_clk;
	wire buf_rdata_clk;
	reg cmdbuf_wr_en;
	wire cmdbuf_rst;
	wire cmdbuf_full;
	wire cmdbuf_vld;
	wire cmdbuf_write;
	wire [1:0] cmdbuf_size;
	wire [7:0] cmdbuf_wstrb;
	wire [31:0] cmdbuf_addr;
	wire [63:0] cmdbuf_wdata;
	localparam [1:0] IDLE = 2'b00;
	localparam [1:0] PEND = 2'b11;
	localparam [1:0] RD = 2'b10;
	localparam [1:0] WR = 2'b01;
	always @(*) begin
		buf_nxtstate = IDLE;
		buf_state_en = 1'b0;
		buf_rdata_en = 1'b0;
		buf_read_error_in = 1'b0;
		cmdbuf_wr_en = 1'b0;
		case (buf_state)
			IDLE: begin
				buf_nxtstate = (ahb_hwrite ? WR : RD);
				buf_state_en = (ahb_hready & ahb_htrans[1]) & ahb_hsel;
			end
			WR: begin
				buf_nxtstate = ((ahb_hresp | (ahb_htrans[1:0] == 2'b00)) | ~ahb_hsel ? IDLE : (ahb_hwrite ? WR : RD));
				buf_state_en = ~cmdbuf_full | ahb_hresp;
				cmdbuf_wr_en = ~cmdbuf_full & ~(ahb_hresp | ((ahb_htrans[1:0] == 2'b01) & ahb_hsel));
			end
			RD: begin
				buf_nxtstate = (ahb_hresp ? IDLE : PEND);
				buf_state_en = ~cmdbuf_full | ahb_hresp;
				cmdbuf_wr_en = ~ahb_hresp & ~cmdbuf_full;
			end
			PEND: begin
				buf_nxtstate = IDLE;
				buf_state_en = axi_rvalid & ~cmdbuf_write;
				buf_rdata_en = buf_state_en;
				buf_read_error_in = buf_state_en & |axi_rresp[1:0];
			end
		endcase
	end
	rvdffs_fpga #(.WIDTH(2)) state_reg(
		.rst_l(rst_l),
		.din(buf_nxtstate),
		.dout({buf_state}),
		.en(buf_state_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk)
	);
	assign master_wstrb[7:0] = ((({8 {ahb_hsize_q[2:0] == 3'b000}} & (8'b00000001 << ahb_haddr_q[2:0])) | ({8 {ahb_hsize_q[2:0] == 3'b001}} & (8'b00000011 << ahb_haddr_q[2:0]))) | ({8 {ahb_hsize_q[2:0] == 3'b010}} & (8'b00001111 << ahb_haddr_q[2:0]))) | ({8 {ahb_hsize_q[2:0] == 3'b011}} & 8'b11111111);
	assign ahb_hreadyout = (ahb_hresp ? ahb_hresp_q & ~ahb_hready_q : ((~cmdbuf_full | (buf_state == IDLE)) & ~((buf_state == RD) | (buf_state == PEND))) & ~buf_read_error);
	assign ahb_hready = ahb_hreadyout & ahb_hreadyin;
	assign ahb_htrans_in[1:0] = {2 {ahb_hsel}} & ahb_htrans[1:0];
	assign ahb_hrdata[63:0] = buf_rdata[63:0];
	assign ahb_hresp = ((((ahb_htrans_q[1:0] != 2'b00) & (buf_state != IDLE)) & ((((~(ahb_addr_in_dccm | ahb_addr_in_iccm) | ((ahb_addr_in_iccm | (ahb_addr_in_dccm & ahb_hwrite_q)) & ~((ahb_hsize_q[1:0] == 2'b10) | (ahb_hsize_q[1:0] == 2'b11)))) | ((ahb_hsize_q[2:0] == 3'h1) & ahb_haddr_q[0])) | ((ahb_hsize_q[2:0] == 3'h2) & |ahb_haddr_q[1:0])) | ((ahb_hsize_q[2:0] == 3'h3) & |ahb_haddr_q[2:0]))) | buf_read_error) | (ahb_hresp_q & ~ahb_hready_q);
	rvdff_fpga #(.WIDTH(64)) buf_rdata_ff(
		.din(axi_rdata[63:0]),
		.dout(buf_rdata[63:0]),
		.clk(buf_rdata_clk),
		.clken(buf_rdata_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) buf_read_error_ff(
		.din(buf_read_error_in),
		.dout(buf_read_error),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hresp_ff(
		.din(ahb_hresp),
		.dout(ahb_hresp_q),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hready_ff(
		.din(ahb_hready),
		.dout(ahb_hready_q),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(2)) htrans_ff(
		.din(ahb_htrans_in[1:0]),
		.dout(ahb_htrans_q[1:0]),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(3)) hsize_ff(
		.din(ahb_hsize[2:0]),
		.dout(ahb_hsize_q[2:0]),
		.clk(ahb_addr_clk),
		.clken(ahb_addr_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hwrite_ff(
		.din(ahb_hwrite),
		.dout(ahb_hwrite_q),
		.clk(ahb_addr_clk),
		.clken(ahb_addr_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(32)) haddr_ff(
		.din(ahb_haddr[31:0]),
		.dout(ahb_haddr_q[31:0]),
		.clk(ahb_addr_clk),
		.clken(ahb_addr_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvrangecheck #(
		.CCM_SADR(pt[1325-:36]),
		.CCM_SIZE(pt[1289-:14])
	) addr_dccm_rangecheck(
		.addr(ahb_haddr_q[31:0]),
		.in_range(ahb_addr_in_dccm),
		.in_region(ahb_addr_in_dccm_region_nc)
	);
	generate
		if (pt[927-:5] == 1) begin : GenICCM
			rvrangecheck #(
				.CCM_SADR(pt[887-:36]),
				.CCM_SIZE(pt[851-:14])
			) addr_iccm_rangecheck(
				.addr(ahb_haddr_q[31:0]),
				.in_range(ahb_addr_in_iccm),
				.in_region(ahb_addr_in_iccm_region_nc)
			);
		end
		else begin : GenNoICCM
			assign ahb_addr_in_iccm = 1'b0;
			assign ahb_addr_in_iccm_region_nc = 1'b0;
		end
	endgenerate
	rvrangecheck #(
		.CCM_SADR(pt[130-:36]),
		.CCM_SIZE(pt[69-:13])
	) addr_pic_rangecheck(
		.addr(ahb_haddr_q[31:0]),
		.in_range(ahb_addr_in_pic),
		.in_region(ahb_addr_in_pic_region_nc)
	);
	assign cmdbuf_rst = (((axi_awvalid & axi_awready) | (axi_arvalid & axi_arready)) & ~cmdbuf_wr_en) | (ahb_hresp & ~cmdbuf_write);
	assign cmdbuf_full = cmdbuf_vld & ~((axi_awvalid & axi_awready) | (axi_arvalid & axi_arready));
	rvdffsc_fpga #(.WIDTH(1)) cmdbuf_vldff(
		.din(1'b1),
		.dout(cmdbuf_vld),
		.en(cmdbuf_wr_en),
		.clear(cmdbuf_rst),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) cmdbuf_writeff(
		.din(ahb_hwrite_q),
		.dout(cmdbuf_write),
		.en(cmdbuf_wr_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(2)) cmdbuf_sizeff(
		.din(ahb_hsize_q[1:0]),
		.dout(cmdbuf_size[1:0]),
		.en(cmdbuf_wr_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(8)) cmdbuf_wstrbff(
		.din(master_wstrb[7:0]),
		.dout(cmdbuf_wstrb[7:0]),
		.en(cmdbuf_wr_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) cmdbuf_addrff(
		.din(ahb_haddr_q[31:0]),
		.dout(cmdbuf_addr[31:0]),
		.en(cmdbuf_wr_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffe #(.WIDTH(64)) cmdbuf_wdataff(
		.din(ahb_hwdata[63:0]),
		.dout(cmdbuf_wdata[63:0]),
		.en(cmdbuf_wr_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	assign axi_awvalid = cmdbuf_vld & cmdbuf_write;
	assign axi_awid[TAG - 1:0] = {TAG {1'sb0}};
	assign axi_awaddr[31:0] = cmdbuf_addr[31:0];
	assign axi_awsize[2:0] = {1'b0, cmdbuf_size[1:0]};
	assign axi_awprot[2:0] = 3'b000;
	assign axi_awlen[7:0] = {8 {1'sb0}};
	assign axi_awburst[1:0] = 2'b01;
	assign axi_wvalid = cmdbuf_vld & cmdbuf_write;
	assign axi_wdata[63:0] = cmdbuf_wdata[63:0];
	assign axi_wstrb[7:0] = cmdbuf_wstrb[7:0];
	assign axi_wlast = 1'b1;
	assign axi_bready = 1'b1;
	assign axi_arvalid = cmdbuf_vld & ~cmdbuf_write;
	assign axi_arid[TAG - 1:0] = {TAG {1'sb0}};
	assign axi_araddr[31:0] = cmdbuf_addr[31:0];
	assign axi_arsize[2:0] = {1'b0, cmdbuf_size[1:0]};
	assign axi_arprot = 3'b000;
	assign axi_arlen[7:0] = {8 {1'sb0}};
	assign axi_arburst[1:0] = 2'b01;
	assign axi_rready = 1'b1;
	assign ahb_addr_clk_en = bus_clk_en & (ahb_hready & ahb_htrans[1]);
	assign buf_rdata_clk_en = bus_clk_en & buf_rdata_en;
	rvclkhdr bus_cgc(
		.en(bus_clk_en),
		.l1clk(bus_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr ahb_addr_cgc(
		.en(ahb_addr_clk_en),
		.l1clk(ahb_addr_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr buf_rdata_cgc(
		.en(buf_rdata_clk_en),
		.l1clk(buf_rdata_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
endmodule
module dmi_jtag_to_core_sync (
	rd_en,
	wr_en,
	rst_n,
	clk,
	reg_en,
	reg_wr_en
);
	input rd_en;
	input wr_en;
	input rst_n;
	input clk;
	output reg_en;
	output reg_wr_en;
	wire c_rd_en;
	wire c_wr_en;
	reg [2:0] rden;
	reg [2:0] wren;
	assign reg_en = c_wr_en | c_rd_en;
	assign reg_wr_en = c_wr_en;
	always @(posedge clk or negedge rst_n)
		if (!rst_n) begin
			rden <= {3 {1'sb0}};
			wren <= {3 {1'sb0}};
		end
		else begin
			rden <= {rden[1:0], rd_en};
			wren <= {wren[1:0], wr_en};
		end
	assign c_rd_en = rden[1] & ~rden[2];
	assign c_wr_en = wren[1] & ~wren[2];
endmodule
module axi4_to_ahb (
	clk,
	free_clk,
	rst_l,
	scan_mode,
	bus_clk_en,
	clk_override,
	dec_tlu_force_halt,
	axi_awvalid,
	axi_awready,
	axi_awid,
	axi_awaddr,
	axi_awsize,
	axi_awprot,
	axi_wvalid,
	axi_wready,
	axi_wdata,
	axi_wstrb,
	axi_wlast,
	axi_bvalid,
	axi_bready,
	axi_bresp,
	axi_bid,
	axi_arvalid,
	axi_arready,
	axi_arid,
	axi_araddr,
	axi_arsize,
	axi_arprot,
	axi_rvalid,
	axi_rready,
	axi_rid,
	axi_rdata,
	axi_rresp,
	axi_rlast,
	ahb_haddr,
	ahb_hburst,
	ahb_hmastlock,
	ahb_hprot,
	ahb_hsize,
	ahb_htrans,
	ahb_hwrite,
	ahb_hwdata,
	ahb_hrdata,
	ahb_hready,
	ahb_hresp
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	parameter TAG = 1;
	input clk;
	input free_clk;
	input rst_l;
	input scan_mode;
	input bus_clk_en;
	input clk_override;
	input dec_tlu_force_halt;
	input wire axi_awvalid;
	output wire axi_awready;
	input wire [TAG - 1:0] axi_awid;
	input wire [31:0] axi_awaddr;
	input wire [2:0] axi_awsize;
	input wire [2:0] axi_awprot;
	input wire axi_wvalid;
	output wire axi_wready;
	input wire [63:0] axi_wdata;
	input wire [7:0] axi_wstrb;
	input wire axi_wlast;
	output wire axi_bvalid;
	input wire axi_bready;
	output wire [1:0] axi_bresp;
	output wire [TAG - 1:0] axi_bid;
	input wire axi_arvalid;
	output wire axi_arready;
	input wire [TAG - 1:0] axi_arid;
	input wire [31:0] axi_araddr;
	input wire [2:0] axi_arsize;
	input wire [2:0] axi_arprot;
	output wire axi_rvalid;
	input wire axi_rready;
	output wire [TAG - 1:0] axi_rid;
	output wire [63:0] axi_rdata;
	output wire [1:0] axi_rresp;
	output wire axi_rlast;
	output wire [31:0] ahb_haddr;
	output wire [2:0] ahb_hburst;
	output wire ahb_hmastlock;
	output wire [3:0] ahb_hprot;
	output wire [2:0] ahb_hsize;
	output reg [1:0] ahb_htrans;
	output wire ahb_hwrite;
	output wire [63:0] ahb_hwdata;
	input wire [63:0] ahb_hrdata;
	input wire ahb_hready;
	input wire ahb_hresp;
	localparam ID = 1;
	localparam PRTY = 1;
	wire [2:0] buf_state;
	reg [2:0] buf_nxtstate;
	wire slave_valid;
	wire slave_ready;
	wire [TAG - 1:0] slave_tag;
	wire [63:0] slave_rdata;
	wire [3:0] slave_opc;
	wire wrbuf_en;
	wire wrbuf_data_en;
	wire wrbuf_cmd_sent;
	wire wrbuf_rst;
	wire wrbuf_vld;
	wire wrbuf_data_vld;
	wire [TAG - 1:0] wrbuf_tag;
	wire [2:0] wrbuf_size;
	wire [31:0] wrbuf_addr;
	wire [63:0] wrbuf_data;
	wire [7:0] wrbuf_byteen;
	wire master_valid;
	reg master_ready;
	wire [TAG - 1:0] master_tag;
	wire [31:0] master_addr;
	wire [63:0] master_wdata;
	wire [2:0] master_size;
	wire [2:0] master_opc;
	wire [7:0] master_byteen;
	wire [31:0] buf_addr;
	wire [1:0] buf_size;
	wire buf_write;
	wire [7:0] buf_byteen;
	wire buf_aligned;
	wire [63:0] buf_data;
	wire [TAG - 1:0] buf_tag;
	wire buf_rst;
	wire [TAG - 1:0] buf_tag_in;
	wire [31:0] buf_addr_in;
	wire [7:0] buf_byteen_in;
	wire [63:0] buf_data_in;
	reg buf_write_in;
	wire buf_aligned_in;
	wire [2:0] buf_size_in;
	reg buf_state_en;
	reg buf_wr_en;
	reg buf_data_wr_en;
	reg slvbuf_error_en;
	wire wr_cmd_vld;
	wire cmd_done_rst;
	reg cmd_done;
	wire cmd_doneQ;
	reg trxn_done;
	reg [2:0] buf_cmd_byte_ptr;
	wire [2:0] buf_cmd_byte_ptrQ;
	wire [2:0] buf_cmd_nxtbyte_ptr;
	reg buf_cmd_byte_ptr_en;
	wire found;
	reg slave_valid_pre;
	wire ahb_hready_q;
	wire ahb_hresp_q;
	wire [1:0] ahb_htrans_q;
	wire ahb_hwrite_q;
	wire [63:0] ahb_hrdata_q;
	wire slvbuf_write;
	wire slvbuf_error;
	wire [TAG - 1:0] slvbuf_tag;
	reg slvbuf_error_in;
	reg slvbuf_wr_en;
	reg bypass_en;
	reg rd_bypass_idle;
	wire last_addr_en;
	wire [31:0] last_bus_addr;
	wire buf_clken;
	wire ahbm_data_clken;
	wire buf_clk;
	wire bus_clk;
	wire ahbm_data_clk;
	wire dec_tlu_force_halt_bus;
	wire dec_tlu_force_halt_bus_ns;
	wire dec_tlu_force_halt_bus_q;
	function automatic [1:0] get_write_size;
		input reg [7:0] byteen;
		reg [1:0] size;
		begin
			size[1:0] = ((2'b11 & {2 {byteen[7:0] == 8'hff}}) | (2'b10 & {2 {(byteen[7:0] == 8'hf0) | (byteen[7:0] == 8'h0f)}})) | (2'b01 & {2 {(((byteen[7:0] == 8'hc0) | (byteen[7:0] == 8'h30)) | (byteen[7:0] == 8'h0c)) | (byteen[7:0] == 8'h03)}});
			get_write_size = size[1:0];
		end
	endfunction
	function automatic [2:0] get_write_addr;
		input reg [7:0] byteen;
		reg [2:0] addr;
		begin
			addr[2:0] = (((3'h0 & {3 {((byteen[7:0] == 8'hff) | (byteen[7:0] == 8'h0f)) | (byteen[7:0] == 8'h03)}}) | (3'h2 & {3 {byteen[7:0] == 8'h0c}})) | (3'h4 & {3 {(byteen[7:0] == 8'hf0) | (byteen[7:0] == 8'h03)}})) | (3'h6 & {3 {byteen[7:0] == 8'hc0}});
			get_write_addr = addr[2:0];
		end
	endfunction
	function automatic signed [2:0] sv2v_cast_3_signed;
		input reg signed [2:0] inp;
		sv2v_cast_3_signed = inp;
	endfunction
	function automatic [2:0] get_nxtbyte_ptr;
		input reg [2:0] current_byte_ptr;
		input reg [7:0] byteen;
		input reg get_next;
		reg [2:0] start_ptr;
		reg found;
		begin
			found = 1'b0;
			start_ptr[2:0] = (get_next ? current_byte_ptr[2:0] + 3'b001 : current_byte_ptr[2:0]);
			begin : sv2v_autoblock_36
				reg signed [31:0] j;
				for (j = 0; j < 8; j = j + 1)
					if (~found) begin
						get_nxtbyte_ptr[2:0] = sv2v_cast_3_signed(j);
						found = found | (byteen[j] & (sv2v_cast_3_signed(j) >= start_ptr[2:0]));
					end
			end
		end
	endfunction
	assign dec_tlu_force_halt_bus = dec_tlu_force_halt | dec_tlu_force_halt_bus_q;
	assign dec_tlu_force_halt_bus_ns = ~bus_clk_en & dec_tlu_force_halt_bus;
	rvdff #(.WIDTH(1)) force_halt_busff(
		.din(dec_tlu_force_halt_bus_ns),
		.dout(dec_tlu_force_halt_bus_q),
		.clk(free_clk),
		.rst_l(rst_l)
	);
	assign wrbuf_en = (axi_awvalid & axi_awready) & master_ready;
	assign wrbuf_data_en = (axi_wvalid & axi_wready) & master_ready;
	assign wrbuf_cmd_sent = (master_valid & master_ready) & (master_opc[2:1] == 2'b01);
	assign wrbuf_rst = (wrbuf_cmd_sent & ~wrbuf_en) | dec_tlu_force_halt_bus;
	assign axi_awready = ~(wrbuf_vld & ~wrbuf_cmd_sent) & master_ready;
	assign axi_wready = ~(wrbuf_data_vld & ~wrbuf_cmd_sent) & master_ready;
	assign axi_arready = ~(wrbuf_vld & wrbuf_data_vld) & master_ready;
	assign axi_rlast = 1'b1;
	assign wr_cmd_vld = wrbuf_vld & wrbuf_data_vld;
	assign master_valid = wr_cmd_vld | axi_arvalid;
	assign master_tag[TAG - 1:0] = (wr_cmd_vld ? wrbuf_tag[TAG - 1:0] : axi_arid[TAG - 1:0]);
	assign master_opc[2:0] = (wr_cmd_vld ? 3'b011 : 3'b000);
	assign master_addr[31:0] = (wr_cmd_vld ? wrbuf_addr[31:0] : axi_araddr[31:0]);
	assign master_size[2:0] = (wr_cmd_vld ? wrbuf_size[2:0] : axi_arsize[2:0]);
	assign master_byteen[7:0] = wrbuf_byteen[7:0];
	assign master_wdata[63:0] = wrbuf_data[63:0];
	assign axi_bvalid = (slave_valid & slave_ready) & slave_opc[3];
	assign axi_bresp[1:0] = (slave_opc[0] ? 2'b10 : (slave_opc[1] ? 2'b11 : 2'b00));
	assign axi_bid[TAG - 1:0] = slave_tag[TAG - 1:0];
	assign axi_rvalid = (slave_valid & slave_ready) & (slave_opc[3:2] == 2'b00);
	assign axi_rresp[1:0] = (slave_opc[0] ? 2'b10 : (slave_opc[1] ? 2'b11 : 2'b00));
	assign axi_rid[TAG - 1:0] = slave_tag[TAG - 1:0];
	assign axi_rdata[63:0] = slave_rdata[63:0];
	assign slave_ready = axi_bready & axi_rready;
	localparam [2:0] CMD_RD = 3'b001;
	localparam [2:0] CMD_WR = 3'b010;
	localparam [2:0] DATA_RD = 3'b011;
	localparam [2:0] DATA_WR = 3'b100;
	localparam [2:0] DONE = 3'b101;
	localparam [2:0] IDLE = 3'b000;
	localparam [2:0] STREAM_ERR_RD = 3'b111;
	localparam [2:0] STREAM_RD = 3'b110;
	always @(*) begin
		buf_nxtstate = IDLE;
		buf_state_en = 1'b0;
		buf_wr_en = 1'b0;
		buf_data_wr_en = 1'b0;
		slvbuf_error_in = 1'b0;
		slvbuf_error_en = 1'b0;
		buf_write_in = 1'b0;
		cmd_done = 1'b0;
		trxn_done = 1'b0;
		buf_cmd_byte_ptr_en = 1'b0;
		buf_cmd_byte_ptr[2:0] = {3 {1'sb0}};
		slave_valid_pre = 1'b0;
		master_ready = 1'b0;
		ahb_htrans[1:0] = 2'b00;
		slvbuf_wr_en = 1'b0;
		bypass_en = 1'b0;
		rd_bypass_idle = 1'b0;
		case (buf_state)
			IDLE: begin
				master_ready = 1'b1;
				buf_write_in = master_opc[2:1] == 2'b01;
				buf_nxtstate = (buf_write_in ? CMD_WR : CMD_RD);
				buf_state_en = master_valid & master_ready;
				buf_wr_en = buf_state_en;
				buf_data_wr_en = buf_state_en & (buf_nxtstate == CMD_WR);
				buf_cmd_byte_ptr_en = buf_state_en;
				buf_cmd_byte_ptr[2:0] = (buf_write_in ? get_nxtbyte_ptr(3'b000, buf_byteen_in[7:0], 1'b0) : master_addr[2:0]);
				bypass_en = buf_state_en;
				rd_bypass_idle = bypass_en & (buf_nxtstate == CMD_RD);
				ahb_htrans[1:0] = {2 {bypass_en}} & 2'b10;
			end
			CMD_RD: begin
				buf_nxtstate = (master_valid & (master_opc[2:0] == 3'b000) ? STREAM_RD : DATA_RD);
				buf_state_en = (ahb_hready_q & (ahb_htrans_q[1:0] != 2'b00)) & ~ahb_hwrite_q;
				cmd_done = buf_state_en & ~master_valid;
				slvbuf_wr_en = buf_state_en;
				master_ready = buf_state_en & (buf_nxtstate == STREAM_RD);
				buf_wr_en = master_ready;
				bypass_en = master_ready & master_valid;
				buf_cmd_byte_ptr[2:0] = (bypass_en ? master_addr[2:0] : buf_addr[2:0]);
				ahb_htrans[1:0] = 2'b10 & {2 {~buf_state_en | bypass_en}};
			end
			STREAM_RD: begin
				master_ready = (ahb_hready_q & ~ahb_hresp_q) & ~(master_valid & (master_opc[2:1] == 2'b01));
				buf_wr_en = (master_valid & master_ready) & (master_opc[2:0] == 3'b000);
				buf_nxtstate = (ahb_hresp_q ? STREAM_ERR_RD : (buf_wr_en ? STREAM_RD : DATA_RD));
				buf_state_en = ahb_hready_q | ahb_hresp_q;
				buf_data_wr_en = buf_state_en;
				slvbuf_error_in = ahb_hresp_q;
				slvbuf_error_en = buf_state_en;
				slave_valid_pre = buf_state_en & ~ahb_hresp_q;
				cmd_done = buf_state_en & ~master_valid;
				bypass_en = ((master_ready & master_valid) & (buf_nxtstate == STREAM_RD)) & buf_state_en;
				buf_cmd_byte_ptr[2:0] = (bypass_en ? master_addr[2:0] : buf_addr[2:0]);
				ahb_htrans[1:0] = 2'b10 & {2 {~((buf_nxtstate != STREAM_RD) & buf_state_en)}};
				slvbuf_wr_en = buf_wr_en;
			end
			STREAM_ERR_RD: begin
				buf_nxtstate = DATA_RD;
				buf_state_en = (ahb_hready_q & (ahb_htrans_q[1:0] != 2'b00)) & ~ahb_hwrite_q;
				slave_valid_pre = buf_state_en;
				slvbuf_wr_en = buf_state_en;
				buf_cmd_byte_ptr[2:0] = buf_addr[2:0];
				ahb_htrans[1:0] = 2'b10 & {2 {~buf_state_en}};
			end
			DATA_RD: begin
				buf_nxtstate = DONE;
				buf_state_en = ahb_hready_q | ahb_hresp_q;
				buf_data_wr_en = buf_state_en;
				slvbuf_error_in = ahb_hresp_q;
				slvbuf_error_en = buf_state_en;
				slvbuf_wr_en = buf_state_en;
			end
			CMD_WR: begin
				buf_nxtstate = DATA_WR;
				trxn_done = (ahb_hready_q & ahb_hwrite_q) & (ahb_htrans_q[1:0] != 2'b00);
				buf_state_en = trxn_done;
				buf_cmd_byte_ptr_en = buf_state_en;
				slvbuf_wr_en = buf_state_en;
				buf_cmd_byte_ptr = (trxn_done ? get_nxtbyte_ptr(buf_cmd_byte_ptrQ[2:0], buf_byteen[7:0], 1'b1) : buf_cmd_byte_ptrQ);
				cmd_done = trxn_done & ((buf_aligned | (buf_cmd_byte_ptrQ == 3'b111)) | (buf_byteen[get_nxtbyte_ptr(buf_cmd_byte_ptrQ[2:0], buf_byteen[7:0], 1'b1)] == 1'b0));
				ahb_htrans[1:0] = {2 {~(cmd_done | cmd_doneQ)}} & 2'b10;
			end
			DATA_WR: begin
				buf_state_en = (cmd_doneQ & ahb_hready_q) | ahb_hresp_q;
				master_ready = (buf_state_en & ~ahb_hresp_q) & slave_ready;
				buf_nxtstate = (ahb_hresp_q | ~slave_ready ? DONE : (master_valid & master_ready ? (master_opc[2:1] == 2'b01 ? CMD_WR : CMD_RD) : IDLE));
				slvbuf_error_in = ahb_hresp_q;
				slvbuf_error_en = buf_state_en;
				buf_write_in = master_opc[2:1] == 2'b01;
				buf_wr_en = buf_state_en & ((buf_nxtstate == CMD_WR) | (buf_nxtstate == CMD_RD));
				buf_data_wr_en = buf_wr_en;
				cmd_done = ahb_hresp_q | ((ahb_hready_q & (ahb_htrans_q[1:0] != 2'b00)) & ((buf_cmd_byte_ptrQ == 3'b111) | (buf_byteen[get_nxtbyte_ptr(buf_cmd_byte_ptrQ[2:0], buf_byteen[7:0], 1'b1)] == 1'b0)));
				bypass_en = (buf_state_en & buf_write_in) & (buf_nxtstate == CMD_WR);
				ahb_htrans[1:0] = {2 {~(cmd_done | cmd_doneQ) | bypass_en}} & 2'b10;
				slave_valid_pre = buf_state_en & (buf_nxtstate != DONE);
				trxn_done = (ahb_hready_q & ahb_hwrite_q) & (ahb_htrans_q[1:0] != 2'b00);
				buf_cmd_byte_ptr_en = trxn_done | bypass_en;
				buf_cmd_byte_ptr = (bypass_en ? get_nxtbyte_ptr(3'b000, buf_byteen_in[7:0], 1'b0) : (trxn_done ? get_nxtbyte_ptr(buf_cmd_byte_ptrQ[2:0], buf_byteen[7:0], 1'b1) : buf_cmd_byte_ptrQ));
			end
			DONE: begin
				buf_nxtstate = IDLE;
				buf_state_en = slave_ready;
				slvbuf_error_en = 1'b1;
				slave_valid_pre = 1'b1;
			end
		endcase
	end
	assign buf_rst = dec_tlu_force_halt_bus;
	assign cmd_done_rst = slave_valid_pre;
	assign buf_addr_in[31:3] = master_addr[31:3];
	assign buf_addr_in[2:0] = (buf_aligned_in & (master_opc[2:1] == 2'b01) ? get_write_addr(master_byteen[7:0]) : master_addr[2:0]);
	assign buf_tag_in[TAG - 1:0] = master_tag[TAG - 1:0];
	assign buf_byteen_in[7:0] = wrbuf_byteen[7:0];
	assign buf_data_in[63:0] = (buf_state == DATA_RD ? ahb_hrdata_q[63:0] : master_wdata[63:0]);
	assign buf_size_in[1:0] = ((buf_aligned_in & (master_size[1:0] == 2'b11)) & (master_opc[2:1] == 2'b01) ? get_write_size(master_byteen[7:0]) : master_size[1:0]);
	assign buf_aligned_in = ((((master_opc[2:0] == 3'b000) | (master_size[1:0] == 2'b00)) | (master_size[1:0] == 2'b01)) | (master_size[1:0] == 2'b10)) | ((master_size[1:0] == 2'b11) & (((((((master_byteen[7:0] == 8'h03) | (master_byteen[7:0] == 8'h0c)) | (master_byteen[7:0] == 8'h30)) | (master_byteen[7:0] == 8'hc0)) | (master_byteen[7:0] == 8'h0f)) | (master_byteen[7:0] == 8'hf0)) | (master_byteen[7:0] == 8'hff)));
	assign ahb_haddr[31:3] = (bypass_en ? master_addr[31:3] : buf_addr[31:3]);
	assign ahb_haddr[2:0] = {3 {ahb_htrans == 2'b10}} & buf_cmd_byte_ptr[2:0];
	assign ahb_hsize[2:0] = (bypass_en ? {1'b0, {2 {buf_aligned_in}} & buf_size_in[1:0]} : {1'b0, {2 {buf_aligned}} & buf_size[1:0]});
	assign ahb_hburst[2:0] = 3'b000;
	assign ahb_hmastlock = 1'b0;
	assign ahb_hprot[3:0] = {3'b001, ~axi_arprot[2]};
	assign ahb_hwrite = (bypass_en ? master_opc[2:1] == 2'b01 : buf_write);
	assign ahb_hwdata[63:0] = buf_data[63:0];
	assign slave_valid = slave_valid_pre;
	assign slave_opc[3:2] = (slvbuf_write ? 2'b11 : 2'b00);
	assign slave_opc[1:0] = {2 {slvbuf_error}} & 2'b10;
	assign slave_rdata[63:0] = (slvbuf_error ? {2 {last_bus_addr[31:0]}} : (buf_state == DONE ? buf_data[63:0] : ahb_hrdata_q[63:0]));
	assign slave_tag[TAG - 1:0] = slvbuf_tag[TAG - 1:0];
	assign last_addr_en = ((ahb_htrans[1:0] != 2'b00) & ahb_hready) & ahb_hwrite;
	rvdffsc_fpga #(.WIDTH(1)) wrbuf_vldff(
		.din(1'b1),
		.dout(wrbuf_vld),
		.en(wrbuf_en),
		.clear(wrbuf_rst),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffsc_fpga #(.WIDTH(1)) wrbuf_data_vldff(
		.din(1'b1),
		.dout(wrbuf_data_vld),
		.en(wrbuf_data_en),
		.clear(wrbuf_rst),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(TAG)) wrbuf_tagff(
		.din(axi_awid[TAG - 1:0]),
		.dout(wrbuf_tag[TAG - 1:0]),
		.en(wrbuf_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(3)) wrbuf_sizeff(
		.din(axi_awsize[2:0]),
		.dout(wrbuf_size[2:0]),
		.en(wrbuf_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) wrbuf_addrff(
		.din(axi_awaddr[31:0]),
		.dout(wrbuf_addr[31:0]),
		.en(wrbuf_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffe #(.WIDTH(64)) wrbuf_dataff(
		.din(axi_wdata[63:0]),
		.dout(wrbuf_data[63:0]),
		.en(wrbuf_data_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffs_fpga #(.WIDTH(8)) wrbuf_byteenff(
		.din(axi_wstrb[7:0]),
		.dout(wrbuf_byteen[7:0]),
		.en(wrbuf_data_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(32)) last_bus_addrff(
		.din(ahb_haddr[31:0]),
		.dout(last_bus_addr[31:0]),
		.en(last_addr_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffsc_fpga #(.WIDTH(3)) buf_state_ff(
		.din(buf_nxtstate),
		.dout({buf_state}),
		.en(buf_state_en),
		.clear(buf_rst),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) buf_writeff(
		.din(buf_write_in),
		.dout(buf_write),
		.en(buf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(TAG)) buf_tagff(
		.din(buf_tag_in[TAG - 1:0]),
		.dout(buf_tag[TAG - 1:0]),
		.en(buf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) buf_addrff(
		.din(buf_addr_in[31:0]),
		.dout(buf_addr[31:0]),
		.en(buf_wr_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffs_fpga #(.WIDTH(2)) buf_sizeff(
		.din(buf_size_in[1:0]),
		.dout(buf_size[1:0]),
		.en(buf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) buf_alignedff(
		.din(buf_aligned_in),
		.dout(buf_aligned),
		.en(buf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(8)) buf_byteenff(
		.din(buf_byteen_in[7:0]),
		.dout(buf_byteen[7:0]),
		.en(buf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(64)) buf_dataff(
		.din(buf_data_in[63:0]),
		.dout(buf_data[63:0]),
		.en(buf_data_wr_en & bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffs_fpga #(.WIDTH(1)) slvbuf_writeff(
		.din(buf_write),
		.dout(slvbuf_write),
		.en(slvbuf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(TAG)) slvbuf_tagff(
		.din(buf_tag[TAG - 1:0]),
		.dout(slvbuf_tag[TAG - 1:0]),
		.en(slvbuf_wr_en),
		.clk(buf_clk),
		.clken(buf_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) slvbuf_errorff(
		.din(slvbuf_error_in),
		.dout(slvbuf_error),
		.en(slvbuf_error_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffsc_fpga #(.WIDTH(1)) buf_cmd_doneff(
		.din(1'b1),
		.dout(cmd_doneQ),
		.en(cmd_done),
		.clear(cmd_done_rst),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(3)) buf_cmd_byte_ptrff(
		.din(buf_cmd_byte_ptr[2:0]),
		.dout(buf_cmd_byte_ptrQ[2:0]),
		.en(buf_cmd_byte_ptr_en),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hready_ff(
		.din(ahb_hready),
		.dout(ahb_hready_q),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(2)) htrans_ff(
		.din(ahb_htrans[1:0]),
		.dout(ahb_htrans_q[1:0]),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hwrite_ff(
		.din(ahb_hwrite),
		.dout(ahb_hwrite_q),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) hresp_ff(
		.din(ahb_hresp),
		.dout(ahb_hresp_q),
		.clk(bus_clk),
		.clken(bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(64)) hrdata_ff(
		.din(ahb_hrdata[63:0]),
		.dout(ahb_hrdata_q[63:0]),
		.clk(ahbm_data_clk),
		.clken(ahbm_data_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	assign buf_clken = bus_clk_en & ((buf_wr_en | slvbuf_wr_en) | clk_override);
	assign ahbm_data_clken = bus_clk_en & ((buf_state != IDLE) | clk_override);
	rvclkhdr bus_cgc(
		.en(bus_clk_en),
		.l1clk(bus_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr buf_cgc(
		.en(buf_clken),
		.l1clk(buf_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr ahbm_data_cgc(
		.en(ahbm_data_clken),
		.l1clk(ahbm_data_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
endmodule
module eb1_dbg (
	dbg_cmd_addr,
	dbg_cmd_wrdata,
	dbg_cmd_valid,
	dbg_cmd_write,
	dbg_cmd_type,
	dbg_cmd_size,
	dbg_core_rst_l,
	core_dbg_rddata,
	core_dbg_cmd_done,
	core_dbg_cmd_fail,
	dbg_dma_bubble,
	dma_dbg_ready,
	dbg_halt_req,
	dbg_resume_req,
	dec_tlu_debug_mode,
	dec_tlu_dbg_halted,
	dec_tlu_mpc_halted_only,
	dec_tlu_resume_ack,
	dmi_reg_en,
	dmi_reg_addr,
	dmi_reg_wr_en,
	dmi_reg_wdata,
	dmi_reg_rdata,
	sb_axi_awvalid,
	sb_axi_awready,
	sb_axi_awid,
	sb_axi_awaddr,
	sb_axi_awregion,
	sb_axi_awlen,
	sb_axi_awsize,
	sb_axi_awburst,
	sb_axi_awlock,
	sb_axi_awcache,
	sb_axi_awprot,
	sb_axi_awqos,
	sb_axi_wvalid,
	sb_axi_wready,
	sb_axi_wdata,
	sb_axi_wstrb,
	sb_axi_wlast,
	sb_axi_bvalid,
	sb_axi_bready,
	sb_axi_bresp,
	sb_axi_arvalid,
	sb_axi_arready,
	sb_axi_arid,
	sb_axi_araddr,
	sb_axi_arregion,
	sb_axi_arlen,
	sb_axi_arsize,
	sb_axi_arburst,
	sb_axi_arlock,
	sb_axi_arcache,
	sb_axi_arprot,
	sb_axi_arqos,
	sb_axi_rvalid,
	sb_axi_rready,
	sb_axi_rdata,
	sb_axi_rresp,
	dbg_bus_clk_en,
	clk,
	rst_l,
	dbg_rst_l,
	clk_override,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	output wire [31:0] dbg_cmd_addr;
	output wire [31:0] dbg_cmd_wrdata;
	output wire dbg_cmd_valid;
	output wire dbg_cmd_write;
	output wire [1:0] dbg_cmd_type;
	output wire [1:0] dbg_cmd_size;
	output wire dbg_core_rst_l;
	input wire [31:0] core_dbg_rddata;
	input wire core_dbg_cmd_done;
	input wire core_dbg_cmd_fail;
	output wire dbg_dma_bubble;
	input wire dma_dbg_ready;
	output reg dbg_halt_req;
	output reg dbg_resume_req;
	input wire dec_tlu_debug_mode;
	input wire dec_tlu_dbg_halted;
	input wire dec_tlu_mpc_halted_only;
	input wire dec_tlu_resume_ack;
	input wire dmi_reg_en;
	input wire [6:0] dmi_reg_addr;
	input wire dmi_reg_wr_en;
	input wire [31:0] dmi_reg_wdata;
	output wire [31:0] dmi_reg_rdata;
	output wire sb_axi_awvalid;
	input wire sb_axi_awready;
	output wire [pt[12-:8] - 1:0] sb_axi_awid;
	output wire [31:0] sb_axi_awaddr;
	output wire [3:0] sb_axi_awregion;
	output wire [7:0] sb_axi_awlen;
	output wire [2:0] sb_axi_awsize;
	output wire [1:0] sb_axi_awburst;
	output wire sb_axi_awlock;
	output wire [3:0] sb_axi_awcache;
	output wire [2:0] sb_axi_awprot;
	output wire [3:0] sb_axi_awqos;
	output wire sb_axi_wvalid;
	input wire sb_axi_wready;
	output wire [63:0] sb_axi_wdata;
	output wire [7:0] sb_axi_wstrb;
	output wire sb_axi_wlast;
	input wire sb_axi_bvalid;
	output wire sb_axi_bready;
	input wire [1:0] sb_axi_bresp;
	output wire sb_axi_arvalid;
	input wire sb_axi_arready;
	output wire [pt[12-:8] - 1:0] sb_axi_arid;
	output wire [31:0] sb_axi_araddr;
	output wire [3:0] sb_axi_arregion;
	output wire [7:0] sb_axi_arlen;
	output wire [2:0] sb_axi_arsize;
	output wire [1:0] sb_axi_arburst;
	output wire sb_axi_arlock;
	output wire [3:0] sb_axi_arcache;
	output wire [2:0] sb_axi_arprot;
	output wire [3:0] sb_axi_arqos;
	input wire sb_axi_rvalid;
	output wire sb_axi_rready;
	input wire [63:0] sb_axi_rdata;
	input wire [1:0] sb_axi_rresp;
	input wire dbg_bus_clk_en;
	input wire clk;
	input wire rst_l;
	input wire dbg_rst_l;
	input wire clk_override;
	input wire scan_mode;
	wire [3:0] dbg_state;
	reg [3:0] dbg_nxtstate;
	reg dbg_state_en;
	wire [31:0] dmstatus_reg;
	wire [31:0] dmcontrol_reg;
	wire [31:0] command_reg;
	wire [31:0] abstractcs_reg;
	wire [31:0] haltsum0_reg;
	wire [31:0] data0_reg;
	wire [31:0] data1_reg;
	wire [31:0] data0_din;
	wire data0_reg_wren;
	wire data0_reg_wren0;
	wire data0_reg_wren1;
	reg data0_reg_wren2;
	wire [31:0] data1_din;
	wire data1_reg_wren;
	wire data1_reg_wren0;
	wire data1_reg_wren1;
	reg abstractcs_busy_wren;
	reg abstractcs_busy_din;
	wire [2:0] abstractcs_error_din;
	wire abstractcs_error_sel0;
	wire abstractcs_error_sel1;
	wire abstractcs_error_seb1;
	wire abstractcs_error_sel3;
	wire abstractcs_error_sel4;
	wire abstractcs_error_sel5;
	wire abstractcs_error_sel6;
	reg dbg_sb_bus_error;
	wire abstractauto_reg_wren;
	wire [1:0] abstractauto_reg;
	wire dmstatus_resumeack_wren;
	wire dmstatus_resumeack_din;
	wire dmstatus_haveresetn_wren;
	wire dmstatus_resumeack;
	wire dmstatus_unavail;
	wire dmstatus_running;
	wire dmstatus_halted;
	wire dmstatus_havereset;
	wire dmstatus_haveresetn;
	wire resumereq;
	wire dmcontrol_wren;
	wire dmcontrol_wren_Q;
	wire execute_command_ns;
	wire execute_command;
	wire command_wren;
	wire command_regno_wren;
	wire command_transfer_din;
	wire command_postexec_din;
	wire [31:0] command_din;
	wire [3:0] dbg_cmd_addr_incr;
	wire [31:0] dbg_cmd_curr_addr;
	wire [31:0] dbg_cmd_next_addr;
	wire [31:0] dmi_reg_rdata_din;
	wire [3:0] sb_state;
	reg [3:0] sb_nxtstate;
	reg sb_state_en;
	wire sbcs_wren;
	reg sbcs_sbbusy_wren;
	reg sbcs_sbbusy_din;
	wire sbcs_sbbusyerror_wren;
	wire sbcs_sbbusyerror_din;
	reg sbcs_sberror_wren;
	reg [2:0] sbcs_sberror_din;
	wire sbcs_unaligned;
	wire sbcs_illegal_size;
	wire [19:15] sbcs_reg_int;
	wire sbdata0_reg_wren0;
	wire sbdata0_reg_wren1;
	wire sbdata0_reg_wren;
	wire [31:0] sbdata0_din;
	wire sbdata1_reg_wren0;
	wire sbdata1_reg_wren1;
	wire sbdata1_reg_wren;
	wire [31:0] sbdata1_din;
	wire sbaddress0_reg_wren0;
	reg sbaddress0_reg_wren1;
	wire sbaddress0_reg_wren;
	wire [31:0] sbaddress0_reg_din;
	wire [3:0] sbaddress0_incr;
	wire sbreadonaddr_access;
	wire sbreadondata_access;
	wire sbdata0wr_access;
	reg sb_abmem_cmd_done_in;
	reg sb_abmem_data_done_in;
	reg sb_abmem_cmd_done_en;
	reg sb_abmem_data_done_en;
	wire sb_abmem_cmd_done;
	wire sb_abmem_data_done;
	wire [31:0] abmem_addr;
	wire abmem_addr_in_dccm_region;
	wire abmem_addr_in_iccm_region;
	wire abmem_addr_in_pic_region;
	wire abmem_addr_core_local;
	wire abmem_addr_external;
	wire sb_cmd_pending;
	wire sb_abmem_cmd_pending;
	wire sb_abmem_cmd_write;
	wire [2:0] sb_abmem_cmd_size;
	wire [31:0] sb_abmem_cmd_addr;
	wire [31:0] sb_abmem_cmd_wdata;
	wire [2:0] sb_cmd_size;
	wire [31:0] sb_cmd_addr;
	wire [63:0] sb_cmd_wdata;
	wire sb_bus_cmd_read;
	wire sb_bus_cmd_write_addr;
	wire sb_bus_cmd_write_data;
	wire sb_bus_rsp_read;
	wire sb_bus_rsp_write;
	wire sb_bus_rsp_error;
	wire [63:0] sb_bus_rdata;
	wire [31:0] sbcs_reg;
	wire [31:0] sbaddress0_reg;
	wire [31:0] sbdata0_reg;
	wire [31:0] sbdata1_reg;
	wire sb_abmem_cmd_arvalid;
	wire sb_abmem_cmd_awvalid;
	wire sb_abmem_cmd_wvalid;
	wire sb_abmem_read_pend;
	wire sb_cmd_awvalid;
	wire sb_cmd_wvalid;
	wire sb_cmd_arvalid;
	wire sb_read_pend;
	wire [31:0] sb_axi_addr;
	wire [63:0] sb_axi_wrdata;
	wire [2:0] sb_axi_size;
	wire dbg_dm_rst_l;
	wire dbg_free_clken;
	wire dbg_free_clk;
	wire sb_free_clken;
	wire sb_free_clk;
	localparam [3:0] IDLE = 4'h0;
	assign dbg_free_clken = (((((((dmi_reg_en | execute_command) | (dbg_state != IDLE)) | dbg_state_en) | dec_tlu_dbg_halted) | dec_tlu_mpc_halted_only) | dec_tlu_debug_mode) | dbg_halt_req) | clk_override;
	localparam [3:0] SBIDLE = 4'h0;
	assign sb_free_clken = (((dmi_reg_en | execute_command) | sb_state_en) | (sb_state != SBIDLE)) | clk_override;
	rvoclkhdr dbg_free_cgc(
		.en(dbg_free_clken),
		.l1clk(dbg_free_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr sb_free_cgc(
		.en(sb_free_clken),
		.l1clk(sb_free_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign dbg_dm_rst_l = dbg_rst_l & (dmcontrol_reg[0] | scan_mode);
	assign dbg_core_rst_l = ~dmcontrol_reg[1] | scan_mode;
	assign sbcs_reg[31:29] = 3'b001;
	assign sbcs_reg[28:23] = {6 {1'sb0}};
	assign sbcs_reg[19:15] = {sbcs_reg_int[19], ~sbcs_reg_int[18], sbcs_reg_int[17:15]};
	assign sbcs_reg[11:5] = 7'h20;
	assign sbcs_reg[4:0] = 5'b01111;
	assign sbcs_wren = (((dmi_reg_addr == 7'h38) & dmi_reg_en) & dmi_reg_wr_en) & (sb_state == SBIDLE);
	assign sbcs_sbbusyerror_wren = (sbcs_wren & dmi_reg_wdata[22]) | ((sbcs_reg[21] & dmi_reg_en) & (((dmi_reg_wr_en & (dmi_reg_addr == 7'h39)) | (dmi_reg_addr == 7'h3c)) | (dmi_reg_addr == 7'h3d)));
	assign sbcs_sbbusyerror_din = ~(sbcs_wren & dmi_reg_wdata[22]);
	rvdffs #(.WIDTH(1)) sbcs_sbbusyerror_reg(
		.din(sbcs_sbbusyerror_din),
		.dout(sbcs_reg[22]),
		.en(sbcs_sbbusyerror_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	rvdffs #(.WIDTH(1)) sbcs_sbbusy_reg(
		.din(sbcs_sbbusy_din),
		.dout(sbcs_reg[21]),
		.en(sbcs_sbbusy_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	rvdffs #(.WIDTH(1)) sbcs_sbreadonaddr_reg(
		.din(dmi_reg_wdata[20]),
		.dout(sbcs_reg[20]),
		.en(sbcs_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	rvdffs #(.WIDTH(5)) sbcs_misc_reg(
		.din({dmi_reg_wdata[19], ~dmi_reg_wdata[18], dmi_reg_wdata[17:15]}),
		.dout(sbcs_reg_int[19:15]),
		.en(sbcs_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	rvdffs #(.WIDTH(3)) sbcs_error_reg(
		.din(sbcs_sberror_din[2:0]),
		.dout(sbcs_reg[14:12]),
		.en(sbcs_sberror_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	assign sbcs_unaligned = (((sbcs_reg[19:17] == 3'b001) & sbaddress0_reg[0]) | ((sbcs_reg[19:17] == 3'b010) & |sbaddress0_reg[1:0])) | ((sbcs_reg[19:17] == 3'b011) & |sbaddress0_reg[2:0]);
	assign sbcs_illegal_size = sbcs_reg[19];
	assign sbaddress0_incr[3:0] = ((({4 {sbcs_reg[19:17] == 3'h0}} & 4'b0001) | ({4 {sbcs_reg[19:17] == 3'h1}} & 4'b0010)) | ({4 {sbcs_reg[19:17] == 3'h2}} & 4'b0100)) | ({4 {sbcs_reg[19:17] == 3'h3}} & 4'b1000);
	assign sbdata0_reg_wren0 = (dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h3c);
	localparam [3:0] RSP_RD = 4'h7;
	assign sbdata0_reg_wren1 = ((sb_state == RSP_RD) & sb_state_en) & ~sbcs_sberror_wren;
	assign sbdata0_reg_wren = sbdata0_reg_wren0 | sbdata0_reg_wren1;
	assign sbdata1_reg_wren0 = (dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h3d);
	assign sbdata1_reg_wren1 = ((sb_state == RSP_RD) & sb_state_en) & ~sbcs_sberror_wren;
	assign sbdata1_reg_wren = sbdata1_reg_wren0 | sbdata1_reg_wren1;
	assign sbdata0_din[31:0] = ({32 {sbdata0_reg_wren0}} & dmi_reg_wdata[31:0]) | ({32 {sbdata0_reg_wren1}} & sb_bus_rdata[31:0]);
	assign sbdata1_din[31:0] = ({32 {sbdata1_reg_wren0}} & dmi_reg_wdata[31:0]) | ({32 {sbdata1_reg_wren1}} & sb_bus_rdata[63:32]);
	rvdffe #(.WIDTH(32)) dbg_sbdata0_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(sbdata0_din[31:0]),
		.dout(sbdata0_reg[31:0]),
		.en(sbdata0_reg_wren),
		.rst_l(dbg_dm_rst_l)
	);
	rvdffe #(.WIDTH(32)) dbg_sbdata1_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(sbdata1_din[31:0]),
		.dout(sbdata1_reg[31:0]),
		.en(sbdata1_reg_wren),
		.rst_l(dbg_dm_rst_l)
	);
	assign sbaddress0_reg_wren0 = (dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h39);
	assign sbaddress0_reg_wren = sbaddress0_reg_wren0 | sbaddress0_reg_wren1;
	assign sbaddress0_reg_din[31:0] = ({32 {sbaddress0_reg_wren0}} & dmi_reg_wdata[31:0]) | ({32 {sbaddress0_reg_wren1}} & (sbaddress0_reg[31:0] + {28'b0000000000000000000000000000, sbaddress0_incr[3:0]}));
	rvdffe #(.WIDTH(32)) dbg_sbaddress0_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(sbaddress0_reg_din[31:0]),
		.dout(sbaddress0_reg[31:0]),
		.en(sbaddress0_reg_wren),
		.rst_l(dbg_dm_rst_l)
	);
	assign sbreadonaddr_access = ((dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h39)) & sbcs_reg[20];
	assign sbreadondata_access = ((dmi_reg_en & ~dmi_reg_wr_en) & (dmi_reg_addr == 7'h3c)) & sbcs_reg[15];
	assign sbdata0wr_access = (dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h3c);
	assign dmcontrol_wren = ((dmi_reg_addr == 7'h10) & dmi_reg_en) & dmi_reg_wr_en;
	assign dmcontrol_reg[29] = 1'b0;
	assign dmcontrol_reg[27:2] = {26 {1'sb0}};
	assign resumereq = (dmcontrol_reg[30] & ~dmcontrol_reg[31]) & dmcontrol_wren_Q;
	rvdffs #(.WIDTH(4)) dmcontrolff(
		.din({dmi_reg_wdata[31:30], dmi_reg_wdata[28], dmi_reg_wdata[1]}),
		.dout({dmcontrol_reg[31:30], dmcontrol_reg[28], dmcontrol_reg[1]}),
		.en(dmcontrol_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	rvdffs #(.WIDTH(1)) dmcontrol_dmactive_ff(
		.din(dmi_reg_wdata[0]),
		.dout(dmcontrol_reg[0]),
		.en(dmcontrol_wren),
		.rst_l(dbg_rst_l),
		.clk(dbg_free_clk)
	);
	rvdff #(.WIDTH(1)) dmcontrol_wrenff(
		.din(dmcontrol_wren),
		.dout(dmcontrol_wren_Q),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	assign dmstatus_reg[31:20] = {12 {1'sb0}};
	assign dmstatus_reg[19:18] = {2 {dmstatus_havereset}};
	assign dmstatus_reg[15:14] = {2 {1'sb0}};
	assign dmstatus_reg[7] = 1'b1;
	assign dmstatus_reg[6:4] = {3 {1'sb0}};
	assign dmstatus_reg[17:16] = {2 {dmstatus_resumeack}};
	assign dmstatus_reg[13:12] = {2 {dmstatus_unavail}};
	assign dmstatus_reg[11:10] = {2 {dmstatus_running}};
	assign dmstatus_reg[9:8] = {2 {dmstatus_halted}};
	assign dmstatus_reg[3:0] = 4'h2;
	localparam [3:0] RESUMING = 4'h9;
	assign dmstatus_resumeack_wren = ((dbg_state == RESUMING) & dec_tlu_resume_ack) | ((dmstatus_resumeack & resumereq) & dmstatus_halted);
	assign dmstatus_resumeack_din = (dbg_state == RESUMING) & dec_tlu_resume_ack;
	assign dmstatus_haveresetn_wren = ((((dmi_reg_addr == 7'h10) & dmi_reg_wdata[28]) & dmi_reg_en) & dmi_reg_wr_en) & dmcontrol_reg[0];
	assign dmstatus_havereset = ~dmstatus_haveresetn;
	assign dmstatus_unavail = dmcontrol_reg[1] | ~rst_l;
	assign dmstatus_running = ~(dmstatus_unavail | dmstatus_halted);
	rvdffs #(.WIDTH(1)) dmstatus_resumeack_reg(
		.din(dmstatus_resumeack_din),
		.dout(dmstatus_resumeack),
		.en(dmstatus_resumeack_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	rvdff #(.WIDTH(1)) dmstatus_halted_reg(
		.din(dec_tlu_dbg_halted & ~dec_tlu_mpc_halted_only),
		.dout(dmstatus_halted),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	rvdffs #(.WIDTH(1)) dmstatus_haveresetn_reg(
		.din(1'b1),
		.dout(dmstatus_haveresetn),
		.en(dmstatus_haveresetn_wren),
		.rst_l(rst_l),
		.clk(dbg_free_clk)
	);
	assign haltsum0_reg[31:1] = {31 {1'sb0}};
	assign haltsum0_reg[0] = dmstatus_halted;
	assign abstractcs_reg[31:13] = {19 {1'sb0}};
	assign abstractcs_reg[11] = 1'b0;
	assign abstractcs_reg[7:4] = {4 {1'sb0}};
	assign abstractcs_reg[3:0] = 4'h2;
	assign abstractcs_error_sel0 = ((abstractcs_reg[12] & ~(|abstractcs_reg[10:8])) & dmi_reg_en) & ((((dmi_reg_wr_en & ((dmi_reg_addr == 7'h16) | (dmi_reg_addr == 7'h17))) | (dmi_reg_addr == 7'h18)) | (dmi_reg_addr == 7'h04)) | (dmi_reg_addr == 7'h05));
	assign abstractcs_error_sel1 = (execute_command & ~(|abstractcs_reg[10:8])) & (((~((command_reg[31:24] == 8'b00000000) | (command_reg[31:24] == 8'h02)) | (((command_reg[22:20] == 3'b011) | command_reg[22]) & (command_reg[31:24] == 8'h02))) | ((command_reg[22:20] != 3'b010) & ((command_reg[31:24] == 8'h00) & command_reg[17]))) | ((command_reg[31:24] == 8'h00) & command_reg[18]));
	assign abstractcs_error_seb1 = ((core_dbg_cmd_done & core_dbg_cmd_fail) | ((execute_command & (command_reg[31:24] == 8'h00)) & (((command_reg[15:12] == 4'h1) & (command_reg[11:5] != 0)) | (command_reg[15:13] != 0)))) & ~(|abstractcs_reg[10:8]);
	localparam [3:0] HALTED = 4'h2;
	assign abstractcs_error_sel3 = (execute_command & (dbg_state != HALTED)) & ~(|abstractcs_reg[10:8]);
	assign abstractcs_error_sel4 = (dbg_sb_bus_error & dbg_bus_clk_en) & ~(|abstractcs_reg[10:8]);
	assign abstractcs_error_sel5 = ((execute_command & (command_reg[31:24] == 8'h02)) & ~(|abstractcs_reg[10:8])) & (((command_reg[22:20] == 3'b001) & data1_reg[0]) | ((command_reg[22:20] == 3'b010) & |data1_reg[1:0]));
	assign abstractcs_error_sel6 = ((dmi_reg_addr == 7'h16) & dmi_reg_en) & dmi_reg_wr_en;
	assign abstractcs_error_din[2:0] = (abstractcs_error_sel0 ? 3'b001 : (abstractcs_error_sel1 ? 3'b010 : (abstractcs_error_seb1 ? 3'b011 : (abstractcs_error_sel3 ? 3'b100 : (abstractcs_error_sel4 ? 3'b101 : (abstractcs_error_sel5 ? 3'b111 : (abstractcs_error_sel6 ? ~dmi_reg_wdata[10:8] & abstractcs_reg[10:8] : abstractcs_reg[10:8])))))));
	rvdffs #(.WIDTH(1)) dmabstractcs_busy_reg(
		.din(abstractcs_busy_din),
		.dout(abstractcs_reg[12]),
		.en(abstractcs_busy_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	rvdff #(.WIDTH(3)) dmabstractcs_error_reg(
		.din(abstractcs_error_din[2:0]),
		.dout(abstractcs_reg[10:8]),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	assign abstractauto_reg_wren = ((dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h18)) & ~abstractcs_reg[12];
	rvdffs #(.WIDTH(2)) dbg_abstractauto_reg(
		.din(dmi_reg_wdata[1:0]),
		.dout(abstractauto_reg[1:0]),
		.en(abstractauto_reg_wren),
		.rst_l(dbg_dm_rst_l),
		.clk(dbg_free_clk)
	);
	assign execute_command_ns = command_wren | ((dmi_reg_en & ~abstractcs_reg[12]) & (((dmi_reg_addr == 7'h04) & abstractauto_reg[0]) | ((dmi_reg_addr == 7'h05) & abstractauto_reg[1])));
	assign command_wren = ((dmi_reg_addr == 7'h17) & dmi_reg_en) & dmi_reg_wr_en;
	localparam [3:0] CMD_DONE = 4'h8;
	assign command_regno_wren = command_wren | ((((command_reg[31:24] == 8'h00) & command_reg[19]) & (dbg_state == CMD_DONE)) & ~(|abstractcs_reg[10:8]));
	assign command_postexec_din = (dmi_reg_wdata[31:24] == 8'h00) & dmi_reg_wdata[18];
	assign command_transfer_din = (dmi_reg_wdata[31:24] == 8'h00) & dmi_reg_wdata[17];
	assign command_din[31:16] = {dmi_reg_wdata[31:24], 1'b0, dmi_reg_wdata[22:19], command_postexec_din, command_transfer_din, dmi_reg_wdata[16]};
	assign command_din[15:0] = (command_wren ? dmi_reg_wdata[15:0] : dbg_cmd_next_addr[15:0]);
	rvdff #(.WIDTH(1)) execute_commandff(
		.din(execute_command_ns),
		.dout(execute_command),
		.clk(dbg_free_clk),
		.rst_l(dbg_dm_rst_l)
	);
	rvdffe #(.WIDTH(16)) dmcommand_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(command_din[31:16]),
		.dout(command_reg[31:16]),
		.en(command_wren),
		.rst_l(dbg_dm_rst_l)
	);
	rvdffe #(.WIDTH(16)) dmcommand_regno_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(command_din[15:0]),
		.dout(command_reg[15:0]),
		.en(command_regno_wren),
		.rst_l(dbg_dm_rst_l)
	);
	assign data0_reg_wren0 = (((dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h04)) & (dbg_state == HALTED)) & ~abstractcs_reg[12];
	localparam [3:0] CORE_CMD_WAIT = 4'h4;
	assign data0_reg_wren1 = (core_dbg_cmd_done & (dbg_state == CORE_CMD_WAIT)) & ~command_reg[16];
	assign data0_reg_wren = (data0_reg_wren0 | data0_reg_wren1) | data0_reg_wren2;
	assign data0_din[31:0] = (({32 {data0_reg_wren0}} & dmi_reg_wdata[31:0]) | ({32 {data0_reg_wren1}} & core_dbg_rddata[31:0])) | ({32 {data0_reg_wren2}} & sb_bus_rdata[31:0]);
	rvdffe #(.WIDTH(32)) dbg_data0_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(data0_din[31:0]),
		.dout(data0_reg[31:0]),
		.en(data0_reg_wren),
		.rst_l(dbg_dm_rst_l)
	);
	assign data1_reg_wren0 = (((dmi_reg_en & dmi_reg_wr_en) & (dmi_reg_addr == 7'h05)) & (dbg_state == HALTED)) & ~abstractcs_reg[12];
	assign data1_reg_wren1 = (((dbg_state == CMD_DONE) & (command_reg[31:24] == 8'h02)) & command_reg[19]) & ~(|abstractcs_reg[10:8]);
	assign data1_reg_wren = data1_reg_wren0 | data1_reg_wren1;
	assign data1_din[31:0] = ({32 {data1_reg_wren0}} & dmi_reg_wdata[31:0]) | ({32 {data1_reg_wren1}} & dbg_cmd_next_addr[31:0]);
	rvdffe #(.WIDTH(32)) dbg_data1_reg(
		.clk(clk),
		.scan_mode(scan_mode),
		.din(data1_din[31:0]),
		.dout(data1_reg[31:0]),
		.en(data1_reg_wren),
		.rst_l(dbg_dm_rst_l)
	);
	rvdffs #(.WIDTH(1)) sb_abmem_cmd_doneff(
		.din(sb_abmem_cmd_done_in),
		.dout(sb_abmem_cmd_done),
		.en(sb_abmem_cmd_done_en),
		.clk(dbg_free_clk),
		.rst_l(dbg_dm_rst_l)
	);
	rvdffs #(.WIDTH(1)) sb_abmem_data_doneff(
		.din(sb_abmem_data_done_in),
		.dout(sb_abmem_data_done),
		.en(sb_abmem_data_done_en),
		.clk(dbg_free_clk),
		.rst_l(dbg_dm_rst_l)
	);
	localparam [3:0] CORE_CMD_START = 4'h3;
	localparam [3:0] HALTING = 4'h1;
	localparam [3:0] SB_CMD_RESP = 4'h7;
	localparam [3:0] SB_CMD_SEND = 4'h6;
	localparam [3:0] SB_CMD_START = 4'h5;
	always @(*) begin
		dbg_nxtstate = IDLE;
		dbg_state_en = 1'b0;
		abstractcs_busy_wren = 1'b0;
		abstractcs_busy_din = 1'b0;
		dbg_halt_req = dmcontrol_wren_Q & dmcontrol_reg[31];
		dbg_resume_req = 1'b0;
		dbg_sb_bus_error = 1'b0;
		data0_reg_wren2 = 1'b0;
		sb_abmem_cmd_done_in = 1'b0;
		sb_abmem_data_done_in = 1'b0;
		sb_abmem_cmd_done_en = 1'b0;
		sb_abmem_data_done_en = 1'b0;
		case (dbg_state)
			IDLE: begin
				dbg_nxtstate = (dmstatus_reg[9] | dec_tlu_mpc_halted_only ? HALTED : HALTING);
				dbg_state_en = (dmcontrol_reg[31] | dmstatus_reg[9]) | dec_tlu_mpc_halted_only;
				dbg_halt_req = dmcontrol_reg[31];
			end
			HALTING: begin
				dbg_nxtstate = HALTED;
				dbg_state_en = dmstatus_reg[9] | dec_tlu_mpc_halted_only;
			end
			HALTED: begin
				dbg_nxtstate = (dmstatus_reg[9] ? (resumereq ? RESUMING : ((command_reg[31:24] == 8'h02) & abmem_addr_external ? SB_CMD_START : CORE_CMD_START)) : (dmcontrol_reg[31] ? HALTING : IDLE));
				dbg_state_en = ((dmstatus_reg[9] & resumereq) | execute_command) | ~(dmstatus_reg[9] | dec_tlu_mpc_halted_only);
				abstractcs_busy_wren = dbg_state_en & ((dbg_nxtstate == CORE_CMD_START) | (dbg_nxtstate == SB_CMD_START));
				abstractcs_busy_din = 1'b1;
				dbg_resume_req = dbg_state_en & (dbg_nxtstate == RESUMING);
			end
			CORE_CMD_START: begin
				dbg_nxtstate = (|abstractcs_reg[10:8] | ((command_reg[31:24] == 8'h00) & ~command_reg[17]) ? CMD_DONE : CORE_CMD_WAIT);
				dbg_state_en = (dbg_cmd_valid | |abstractcs_reg[10:8]) | ((command_reg[31:24] == 8'h00) & ~command_reg[17]);
			end
			CORE_CMD_WAIT: begin
				dbg_nxtstate = CMD_DONE;
				dbg_state_en = core_dbg_cmd_done;
			end
			SB_CMD_START: begin
				dbg_nxtstate = (|abstractcs_reg[10:8] ? CMD_DONE : SB_CMD_SEND);
				dbg_state_en = (dbg_bus_clk_en & ~sb_cmd_pending) | |abstractcs_reg[10:8];
			end
			SB_CMD_SEND: begin
				sb_abmem_cmd_done_in = 1'b1;
				sb_abmem_data_done_in = 1'b1;
				sb_abmem_cmd_done_en = (sb_bus_cmd_read | sb_bus_cmd_write_addr) & dbg_bus_clk_en;
				sb_abmem_data_done_en = (sb_bus_cmd_read | sb_bus_cmd_write_data) & dbg_bus_clk_en;
				dbg_nxtstate = SB_CMD_RESP;
				dbg_state_en = ((sb_abmem_cmd_done | sb_abmem_cmd_done_en) & (sb_abmem_data_done | sb_abmem_data_done_en)) & dbg_bus_clk_en;
			end
			SB_CMD_RESP: begin
				dbg_nxtstate = CMD_DONE;
				dbg_state_en = (sb_bus_rsp_read | sb_bus_rsp_write) & dbg_bus_clk_en;
				dbg_sb_bus_error = ((sb_bus_rsp_read | sb_bus_rsp_write) & sb_bus_rsp_error) & dbg_bus_clk_en;
				data0_reg_wren2 = (dbg_state_en & ~sb_abmem_cmd_write) & ~dbg_sb_bus_error;
			end
			CMD_DONE: begin
				dbg_nxtstate = HALTED;
				dbg_state_en = 1'b1;
				abstractcs_busy_wren = dbg_state_en;
				abstractcs_busy_din = 1'b0;
				sb_abmem_cmd_done_in = 1'b0;
				sb_abmem_data_done_in = 1'b0;
				sb_abmem_cmd_done_en = 1'b1;
				sb_abmem_data_done_en = 1'b1;
			end
			RESUMING: begin
				dbg_nxtstate = IDLE;
				dbg_state_en = dmstatus_reg[17];
			end
			default: begin
				dbg_nxtstate = IDLE;
				dbg_state_en = 1'b0;
				abstractcs_busy_wren = 1'b0;
				abstractcs_busy_din = 1'b0;
				dbg_halt_req = 1'b0;
				dbg_resume_req = 1'b0;
				dbg_sb_bus_error = 1'b0;
				data0_reg_wren2 = 1'b0;
				sb_abmem_cmd_done_in = 1'b0;
				sb_abmem_data_done_in = 1'b0;
				sb_abmem_cmd_done_en = 1'b0;
				sb_abmem_data_done_en = 1'b0;
			end
		endcase
	end
	assign dmi_reg_rdata_din[31:0] = ((((((((((({32 {dmi_reg_addr == 7'h04}} & data0_reg[31:0]) | ({32 {dmi_reg_addr == 7'h05}} & data1_reg[31:0])) | ({32 {dmi_reg_addr == 7'h10}} & {2'b00, dmcontrol_reg[29], 1'b0, dmcontrol_reg[27:0]})) | ({32 {dmi_reg_addr == 7'h11}} & dmstatus_reg[31:0])) | ({32 {dmi_reg_addr == 7'h16}} & abstractcs_reg[31:0])) | ({32 {dmi_reg_addr == 7'h17}} & command_reg[31:0])) | ({32 {dmi_reg_addr == 7'h18}} & {30'h00000000, abstractauto_reg[1:0]})) | ({32 {dmi_reg_addr == 7'h40}} & haltsum0_reg[31:0])) | ({32 {dmi_reg_addr == 7'h38}} & sbcs_reg[31:0])) | ({32 {dmi_reg_addr == 7'h39}} & sbaddress0_reg[31:0])) | ({32 {dmi_reg_addr == 7'h3c}} & sbdata0_reg[31:0])) | ({32 {dmi_reg_addr == 7'h3d}} & sbdata1_reg[31:0]);
	rvdffs #(.WIDTH(4)) dbg_state_reg(
		.din(dbg_nxtstate),
		.dout({dbg_state}),
		.en(dbg_state_en),
		.rst_l(dbg_dm_rst_l & rst_l),
		.clk(dbg_free_clk)
	);
	rvdffe #(.WIDTH(32)) dmi_rddata_reg(
		.din(dmi_reg_rdata_din[31:0]),
		.dout(dmi_reg_rdata[31:0]),
		.en(dmi_reg_en),
		.rst_l(dbg_dm_rst_l),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign abmem_addr[31:0] = data1_reg[31:0];
	assign abmem_addr_core_local = (abmem_addr_in_dccm_region | abmem_addr_in_iccm_region) | abmem_addr_in_pic_region;
	assign abmem_addr_external = ~abmem_addr_core_local;
	assign abmem_addr_in_dccm_region = (abmem_addr[31:28] == pt[1333-:8]) & pt[1365-:5];
	assign abmem_addr_in_iccm_region = (abmem_addr[31:28] == pt[895-:8]) & pt[927-:5];
	assign abmem_addr_in_pic_region = abmem_addr[31:28] == pt[77-:8];
	assign dbg_cmd_addr[31:0] = (command_reg[31:24] == 8'h02 ? data1_reg[31:0] : {20'b00000000000000000000, command_reg[11:0]});
	assign dbg_cmd_wrdata[31:0] = data0_reg[31:0];
	assign dbg_cmd_valid = ((dbg_state == CORE_CMD_START) & ~((|abstractcs_reg[10:8] | ((command_reg[31:24] == 8'h00) & ~command_reg[17])) | ((command_reg[31:24] == 8'h02) & abmem_addr_external))) & dma_dbg_ready;
	assign dbg_cmd_write = command_reg[16];
	assign dbg_cmd_type[1:0] = (command_reg[31:24] == 8'h02 ? 2'b10 : {1'b0, command_reg[15:12] == 4'b0000});
	assign dbg_cmd_size[1:0] = command_reg[21:20];
	assign dbg_cmd_addr_incr[3:0] = (command_reg[31:24] == 8'h02 ? 4'h1 << sb_abmem_cmd_size[1:0] : 4'h1);
	assign dbg_cmd_curr_addr[31:0] = (command_reg[31:24] == 8'h02 ? data1_reg[31:0] : {16'b0000000000000000, command_reg[15:0]});
	assign dbg_cmd_next_addr[31:0] = dbg_cmd_curr_addr[31:0] + {28'h0000000, dbg_cmd_addr_incr[3:0]};
	assign dbg_dma_bubble = ((dbg_state == CORE_CMD_START) & ~(|abstractcs_reg[10:8])) | (dbg_state == CORE_CMD_WAIT);
	localparam [3:0] CMD_RD = 4'h3;
	localparam [3:0] CMD_WR = 4'h4;
	localparam [3:0] CMD_WR_ADDR = 4'h5;
	localparam [3:0] CMD_WR_DATA = 4'h6;
	localparam [3:0] RSP_WR = 4'h8;
	assign sb_cmd_pending = (((((sb_state == CMD_RD) | (sb_state == CMD_WR)) | (sb_state == CMD_WR_ADDR)) | (sb_state == CMD_WR_DATA)) | (sb_state == RSP_RD)) | (sb_state == RSP_WR);
	assign sb_abmem_cmd_pending = ((dbg_state == SB_CMD_START) | (dbg_state == SB_CMD_SEND)) | (dbg_state == SB_CMD_RESP);
	localparam [3:0] DONE = 4'h9;
	localparam [3:0] WAIT_RD = 4'h1;
	localparam [3:0] WAIT_WR = 4'h2;
	always @(*) begin
		sb_nxtstate = SBIDLE;
		sb_state_en = 1'b0;
		sbcs_sbbusy_wren = 1'b0;
		sbcs_sbbusy_din = 1'b0;
		sbcs_sberror_wren = 1'b0;
		sbcs_sberror_din[2:0] = 3'b000;
		sbaddress0_reg_wren1 = 1'b0;
		case (sb_state)
			SBIDLE: begin
				sb_nxtstate = (sbdata0wr_access ? WAIT_WR : WAIT_RD);
				sb_state_en = (((sbdata0wr_access | sbreadondata_access) | sbreadonaddr_access) & ~(|sbcs_reg[14:12])) & ~sbcs_reg[22];
				sbcs_sbbusy_wren = sb_state_en;
				sbcs_sbbusy_din = 1'b1;
				sbcs_sberror_wren = sbcs_wren & |dmi_reg_wdata[14:12];
				sbcs_sberror_din[2:0] = ~dmi_reg_wdata[14:12] & sbcs_reg[14:12];
			end
			WAIT_RD: begin
				sb_nxtstate = (sbcs_unaligned | sbcs_illegal_size ? DONE : CMD_RD);
				sb_state_en = ((dbg_bus_clk_en & ~sb_abmem_cmd_pending) | sbcs_unaligned) | sbcs_illegal_size;
				sbcs_sberror_wren = sbcs_unaligned | sbcs_illegal_size;
				sbcs_sberror_din[2:0] = (sbcs_unaligned ? 3'b011 : 3'b100);
			end
			WAIT_WR: begin
				sb_nxtstate = (sbcs_unaligned | sbcs_illegal_size ? DONE : CMD_WR);
				sb_state_en = ((dbg_bus_clk_en & ~sb_abmem_cmd_pending) | sbcs_unaligned) | sbcs_illegal_size;
				sbcs_sberror_wren = sbcs_unaligned | sbcs_illegal_size;
				sbcs_sberror_din[2:0] = (sbcs_unaligned ? 3'b011 : 3'b100);
			end
			CMD_RD: begin
				sb_nxtstate = RSP_RD;
				sb_state_en = sb_bus_cmd_read & dbg_bus_clk_en;
			end
			CMD_WR: begin
				sb_nxtstate = (sb_bus_cmd_write_addr & sb_bus_cmd_write_data ? RSP_WR : (sb_bus_cmd_write_data ? CMD_WR_ADDR : CMD_WR_DATA));
				sb_state_en = (sb_bus_cmd_write_addr | sb_bus_cmd_write_data) & dbg_bus_clk_en;
			end
			CMD_WR_ADDR: begin
				sb_nxtstate = RSP_WR;
				sb_state_en = sb_bus_cmd_write_addr & dbg_bus_clk_en;
			end
			CMD_WR_DATA: begin
				sb_nxtstate = RSP_WR;
				sb_state_en = sb_bus_cmd_write_data & dbg_bus_clk_en;
			end
			RSP_RD: begin
				sb_nxtstate = DONE;
				sb_state_en = sb_bus_rsp_read & dbg_bus_clk_en;
				sbcs_sberror_wren = sb_state_en & sb_bus_rsp_error;
				sbcs_sberror_din[2:0] = 3'b010;
			end
			RSP_WR: begin
				sb_nxtstate = DONE;
				sb_state_en = sb_bus_rsp_write & dbg_bus_clk_en;
				sbcs_sberror_wren = sb_state_en & sb_bus_rsp_error;
				sbcs_sberror_din[2:0] = 3'b010;
			end
			DONE: begin
				sb_nxtstate = SBIDLE;
				sb_state_en = 1'b1;
				sbcs_sbbusy_wren = 1'b1;
				sbcs_sbbusy_din = 1'b0;
				sbaddress0_reg_wren1 = sbcs_reg[16] & (sbcs_reg[14:12] == 3'b000);
			end
			default: begin
				sb_nxtstate = SBIDLE;
				sb_state_en = 1'b0;
				sbcs_sbbusy_wren = 1'b0;
				sbcs_sbbusy_din = 1'b0;
				sbcs_sberror_wren = 1'b0;
				sbcs_sberror_din[2:0] = 3'b000;
				sbaddress0_reg_wren1 = 1'b0;
			end
		endcase
	end
	rvdffs #(.WIDTH(4)) sb_state_reg(
		.din(sb_nxtstate),
		.dout({sb_state}),
		.en(sb_state_en),
		.rst_l(dbg_dm_rst_l),
		.clk(sb_free_clk)
	);
	assign sb_abmem_cmd_write = command_reg[16];
	assign sb_abmem_cmd_size[2:0] = {1'b0, command_reg[21:20]};
	assign sb_abmem_cmd_addr[31:0] = abmem_addr[31:0];
	assign sb_abmem_cmd_wdata[31:0] = data0_reg[31:0];
	assign sb_cmd_size[2:0] = sbcs_reg[19:17];
	assign sb_cmd_wdata[63:0] = {sbdata1_reg[31:0], sbdata0_reg[31:0]};
	assign sb_cmd_addr[31:0] = sbaddress0_reg[31:0];
	assign sb_abmem_cmd_awvalid = ((dbg_state == SB_CMD_SEND) & sb_abmem_cmd_write) & ~sb_abmem_cmd_done;
	assign sb_abmem_cmd_wvalid = ((dbg_state == SB_CMD_SEND) & sb_abmem_cmd_write) & ~sb_abmem_data_done;
	assign sb_abmem_cmd_arvalid = (((dbg_state == SB_CMD_SEND) & ~sb_abmem_cmd_write) & ~sb_abmem_cmd_done) & ~sb_abmem_data_done;
	assign sb_abmem_read_pend = (dbg_state == SB_CMD_RESP) & ~sb_abmem_cmd_write;
	assign sb_cmd_awvalid = (sb_state == CMD_WR) | (sb_state == CMD_WR_ADDR);
	assign sb_cmd_wvalid = (sb_state == CMD_WR) | (sb_state == CMD_WR_DATA);
	assign sb_cmd_arvalid = sb_state == CMD_RD;
	assign sb_read_pend = sb_state == RSP_RD;
	assign sb_axi_size[2:0] = (((sb_abmem_cmd_awvalid | sb_abmem_cmd_wvalid) | sb_abmem_cmd_arvalid) | sb_abmem_read_pend ? sb_abmem_cmd_size[2:0] : sb_cmd_size[2:0]);
	assign sb_axi_addr[31:0] = (((sb_abmem_cmd_awvalid | sb_abmem_cmd_wvalid) | sb_abmem_cmd_arvalid) | sb_abmem_read_pend ? sb_abmem_cmd_addr[31:0] : sb_cmd_addr[31:0]);
	assign sb_axi_wrdata[63:0] = (sb_abmem_cmd_awvalid | sb_abmem_cmd_wvalid ? {2 {sb_abmem_cmd_wdata[31:0]}} : sb_cmd_wdata[63:0]);
	assign sb_bus_cmd_read = sb_axi_arvalid & sb_axi_arready;
	assign sb_bus_cmd_write_addr = sb_axi_awvalid & sb_axi_awready;
	assign sb_bus_cmd_write_data = sb_axi_wvalid & sb_axi_wready;
	assign sb_bus_rsp_read = sb_axi_rvalid & sb_axi_rready;
	assign sb_bus_rsp_write = sb_axi_bvalid & sb_axi_bready;
	assign sb_bus_rsp_error = (sb_bus_rsp_read & |sb_axi_rresp[1:0]) | (sb_bus_rsp_write & |sb_axi_bresp[1:0]);
	assign sb_axi_awvalid = sb_abmem_cmd_awvalid | sb_cmd_awvalid;
	assign sb_axi_awaddr[31:0] = sb_axi_addr[31:0];
	assign sb_axi_awid[pt[12-:8] - 1:0] = {pt[12-:8] {1'sb0}};
	assign sb_axi_awsize[2:0] = sb_axi_size[2:0];
	assign sb_axi_awprot[2:0] = 3'b001;
	assign sb_axi_awcache[3:0] = 4'b1111;
	assign sb_axi_awregion[3:0] = sb_axi_addr[31:28];
	assign sb_axi_awlen[7:0] = {8 {1'sb0}};
	assign sb_axi_awburst[1:0] = 2'b01;
	assign sb_axi_awqos[3:0] = {4 {1'sb0}};
	assign sb_axi_awlock = 1'b0;
	assign sb_axi_wvalid = sb_abmem_cmd_wvalid | sb_cmd_wvalid;
	assign sb_axi_wdata[63:0] = ((({64 {sb_axi_size[2:0] == 3'h0}} & {8 {sb_axi_wrdata[7:0]}}) | ({64 {sb_axi_size[2:0] == 3'h1}} & {4 {sb_axi_wrdata[15:0]}})) | ({64 {sb_axi_size[2:0] == 3'h2}} & {2 {sb_axi_wrdata[31:0]}})) | ({64 {sb_axi_size[2:0] == 3'h3}} & {sb_axi_wrdata[63:0]});
	assign sb_axi_wstrb[7:0] = ((({8 {sb_axi_size[2:0] == 3'h0}} & (8'h01 << sb_axi_addr[2:0])) | ({8 {sb_axi_size[2:0] == 3'h1}} & (8'h03 << {sb_axi_addr[2:1], 1'b0}))) | ({8 {sb_axi_size[2:0] == 3'h2}} & (8'h0f << {sb_axi_addr[2], 2'b00}))) | ({8 {sb_axi_size[2:0] == 3'h3}} & 8'hff);
	assign sb_axi_wlast = 1'b1;
	assign sb_axi_arvalid = sb_abmem_cmd_arvalid | sb_cmd_arvalid;
	assign sb_axi_araddr[31:0] = sb_axi_addr[31:0];
	assign sb_axi_arid[pt[12-:8] - 1:0] = {pt[12-:8] {1'sb0}};
	assign sb_axi_arsize[2:0] = sb_axi_size[2:0];
	assign sb_axi_arprot[2:0] = 3'b001;
	assign sb_axi_arcache[3:0] = 4'b0000;
	assign sb_axi_arregion[3:0] = sb_axi_addr[31:28];
	assign sb_axi_arlen[7:0] = {8 {1'sb0}};
	assign sb_axi_arburst[1:0] = 2'b01;
	assign sb_axi_arqos[3:0] = {4 {1'sb0}};
	assign sb_axi_arlock = 1'b0;
	assign sb_axi_bready = 1'b1;
	assign sb_axi_rready = 1'b1;
	assign sb_bus_rdata[63:0] = ((({64 {sb_axi_size == 3'h0}} & ((sb_axi_rdata[63:0] >> (8 * sb_axi_addr[2:0])) & 64'h00000000000000ff)) | ({64 {sb_axi_size == 3'h1}} & ((sb_axi_rdata[63:0] >> (16 * sb_axi_addr[2:1])) & 64'h000000000000ffff))) | ({64 {sb_axi_size == 3'h2}} & ((sb_axi_rdata[63:0] >> (32 * sb_axi_addr[2])) & 64'h00000000ffffffff))) | ({64 {sb_axi_size == 3'h3}} & sb_axi_rdata[63:0]);
endmodule
module eb1_dec (
	clk,
	active_clk,
	free_clk,
	free_l2clk,
	lsu_fastint_stall_any,
	dec_extint_stall,
	dec_i0_decode_d,
	dec_pause_state_cg,
	dec_tlu_core_empty,
	rst_l,
	rst_vec,
	nmi_int,
	nmi_vec,
	i_cpu_halt_req,
	i_cpu_run_req,
	o_cpu_halt_status,
	o_cpu_halt_ack,
	o_cpu_run_ack,
	o_debug_mode_status,
	core_id,
	mpc_debug_halt_req,
	mpc_debug_run_req,
	mpc_reset_run_req,
	mpc_debug_halt_ack,
	mpc_debug_run_ack,
	debug_brkpt_status,
	exu_pmu_i0_br_misp,
	exu_pmu_i0_br_ataken,
	exu_pmu_i0_pc4,
	lsu_nonblock_load_valid_m,
	lsu_nonblock_load_tag_m,
	lsu_nonblock_load_inv_r,
	lsu_nonblock_load_inv_tag_r,
	lsu_nonblock_load_data_valid,
	lsu_nonblock_load_data_error,
	lsu_nonblock_load_data_tag,
	lsu_nonblock_load_data,
	lsu_pmu_bus_trxn,
	lsu_pmu_bus_misaligned,
	lsu_pmu_bus_error,
	lsu_pmu_bus_busy,
	lsu_pmu_misaligned_m,
	lsu_pmu_load_external_m,
	lsu_pmu_store_external_m,
	dma_pmu_dccm_read,
	dma_pmu_dccm_write,
	dma_pmu_any_read,
	dma_pmu_any_write,
	lsu_fir_addr,
	lsu_fir_error,
	ifu_pmu_instr_aligned,
	ifu_pmu_fetch_stall,
	ifu_pmu_ic_miss,
	ifu_pmu_ic_hit,
	ifu_pmu_bus_error,
	ifu_pmu_bus_busy,
	ifu_pmu_bus_trxn,
	ifu_ic_error_start,
	ifu_iccm_rd_ecc_single_err,
	lsu_trigger_match_m,
	dbg_cmd_valid,
	dbg_cmd_write,
	dbg_cmd_type,
	dbg_cmd_addr,
	dbg_cmd_wrdata,
	ifu_i0_icaf,
	ifu_i0_icaf_type,
	ifu_i0_icaf_second,
	ifu_i0_dbecc,
	lsu_idle_any,
	i0_brp,
	ifu_i0_bp_index,
	ifu_i0_bp_fghr,
	ifu_i0_bp_btag,
	ifu_i0_fa_index,
	lsu_error_pkt_r,
	lsu_single_ecc_error_incr,
	lsu_imprecise_error_load_any,
	lsu_imprecise_error_store_any,
	lsu_imprecise_error_addr_any,
	exu_div_result,
	exu_div_wren,
	exu_csr_rs1_x,
	lsu_result_m,
	lsu_result_corr_r,
	lsu_load_stall_any,
	lsu_store_stall_any,
	dma_dccm_stall_any,
	dma_iccm_stall_any,
	iccm_dma_sb_error,
	exu_flush_final,
	exu_npc_r,
	exu_i0_result_x,
	ifu_i0_valid,
	ifu_i0_instr,
	ifu_i0_pc,
	ifu_i0_pc4,
	exu_i0_pc_x,
	mexintpend,
	timer_int,
	soft_int,
	pic_claimid,
	pic_pl,
	mhwakeup,
	dec_tlu_meicurpl,
	dec_tlu_meipt,
	ifu_ic_debug_rd_data,
	ifu_ic_debug_rd_data_valid,
	dec_tlu_ic_diag_pkt,
	dbg_halt_req,
	dbg_resume_req,
	ifu_miss_state_idle,
	dec_tlu_dbg_halted,
	dec_tlu_debug_mode,
	dec_tlu_resume_ack,
	dec_tlu_flush_noredir_r,
	dec_tlu_mpc_halted_only,
	dec_tlu_flush_leak_one_r,
	dec_tlu_flush_err_r,
	dec_tlu_meihap,
	dec_debug_wdata_rs1_d,
	dec_dbg_rddata,
	dec_dbg_cmd_done,
	dec_dbg_cmd_fail,
	trigger_pkt_any,
	dec_tlu_force_halt,
	exu_i0_br_hist_r,
	exu_i0_br_error_r,
	exu_i0_br_start_error_r,
	exu_i0_br_valid_r,
	exu_i0_br_mp_r,
	exu_i0_br_middle_r,
	exu_i0_br_way_r,
	dec_i0_rs1_en_d,
	dec_i0_rs2_en_d,
	gpr_i0_rs1_d,
	gpr_i0_rs2_d,
	dec_i0_immed_d,
	dec_i0_br_immed_d,
	i0_ap,
	dec_i0_alu_decode_d,
	dec_i0_branch_d,
	dec_i0_select_pc_d,
	dec_i0_pc_d,
	dec_i0_rs1_bypass_en_d,
	dec_i0_rs2_bypass_en_d,
	dec_i0_result_r,
	lsu_p,
	dec_qual_lsu_d,
	mul_p,
	div_p,
	dec_div_cancel,
	dec_lsu_offset_d,
	dec_csr_ren_d,
	dec_csr_rddata_d,
	dec_tlu_flush_lower_r,
	dec_tlu_flush_lower_wb,
	dec_tlu_flush_path_r,
	dec_tlu_i0_kill_writeb_r,
	dec_tlu_fence_i_r,
	pred_correct_npc_x,
	dec_tlu_br0_r_pkt,
	dec_tlu_perfcnt0,
	dec_tlu_perfcnt1,
	dec_tlu_perfcnt2,
	dec_tlu_perfcnt3,
	dec_i0_predict_p_d,
	i0_predict_fghr_d,
	i0_predict_index_d,
	i0_predict_btag_d,
	dec_fa_error_index,
	dec_lsu_valid_raw_d,
	dec_tlu_mrac_ff,
	dec_data_en,
	dec_ctl_en,
	ifu_i0_cinst,
	trace_rv_trace_pkt,
	dec_tlu_external_ldfwd_disable,
	dec_tlu_sideeffect_posted_disable,
	dec_tlu_core_ecc_disable,
	dec_tlu_bpred_disable,
	dec_tlu_wb_coalescing_disable,
	dec_tlu_dma_qos_prty,
	dec_tlu_misc_clk_override,
	dec_tlu_ifu_clk_override,
	dec_tlu_lsu_clk_override,
	dec_tlu_bus_clk_override,
	dec_tlu_pic_clk_override,
	dec_tlu_picio_clk_override,
	dec_tlu_dccm_clk_override,
	dec_tlu_icm_clk_override,
	dec_tlu_i0_commit_cmt,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire active_clk;
	input wire free_clk;
	input wire free_l2clk;
	input wire lsu_fastint_stall_any;
	output wire dec_extint_stall;
	output wire dec_i0_decode_d;
	output wire dec_pause_state_cg;
	output wire dec_tlu_core_empty;
	input wire rst_l;
	input wire [31:1] rst_vec;
	input wire nmi_int;
	input wire [31:1] nmi_vec;
	input wire i_cpu_halt_req;
	input wire i_cpu_run_req;
	output wire o_cpu_halt_status;
	output wire o_cpu_halt_ack;
	output wire o_cpu_run_ack;
	output wire o_debug_mode_status;
	input wire [31:4] core_id;
	input wire mpc_debug_halt_req;
	input wire mpc_debug_run_req;
	input wire mpc_reset_run_req;
	output wire mpc_debug_halt_ack;
	output wire mpc_debug_run_ack;
	output wire debug_brkpt_status;
	input wire exu_pmu_i0_br_misp;
	input wire exu_pmu_i0_br_ataken;
	input wire exu_pmu_i0_pc4;
	input wire lsu_nonblock_load_valid_m;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	input wire lsu_nonblock_load_inv_r;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	input wire lsu_nonblock_load_data_valid;
	input wire lsu_nonblock_load_data_error;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	input wire [31:0] lsu_nonblock_load_data;
	input wire lsu_pmu_bus_trxn;
	input wire lsu_pmu_bus_misaligned;
	input wire lsu_pmu_bus_error;
	input wire lsu_pmu_bus_busy;
	input wire lsu_pmu_misaligned_m;
	input wire lsu_pmu_load_external_m;
	input wire lsu_pmu_store_external_m;
	input wire dma_pmu_dccm_read;
	input wire dma_pmu_dccm_write;
	input wire dma_pmu_any_read;
	input wire dma_pmu_any_write;
	input wire [31:1] lsu_fir_addr;
	input wire [1:0] lsu_fir_error;
	input wire ifu_pmu_instr_aligned;
	input wire ifu_pmu_fetch_stall;
	input wire ifu_pmu_ic_miss;
	input wire ifu_pmu_ic_hit;
	input wire ifu_pmu_bus_error;
	input wire ifu_pmu_bus_busy;
	input wire ifu_pmu_bus_trxn;
	input wire ifu_ic_error_start;
	input wire ifu_iccm_rd_ecc_single_err;
	input wire [3:0] lsu_trigger_match_m;
	input wire dbg_cmd_valid;
	input wire dbg_cmd_write;
	input wire [1:0] dbg_cmd_type;
	input wire [31:0] dbg_cmd_addr;
	input wire [1:0] dbg_cmd_wrdata;
	input wire ifu_i0_icaf;
	input wire [1:0] ifu_i0_icaf_type;
	input wire ifu_i0_icaf_second;
	input wire ifu_i0_dbecc;
	input wire lsu_idle_any;
	input wire [50:0] i0_brp;
	input wire [pt[2172-:9]:pt[2163-:6]] ifu_i0_bp_index;
	input wire [pt[2236-:8] - 1:0] ifu_i0_bp_fghr;
	input wire [pt[2139-:9] - 1:0] ifu_i0_bp_btag;
	input wire [$clog2(pt[2061-:14]) - 1:0] ifu_i0_fa_index;
	input wire [39:0] lsu_error_pkt_r;
	input wire lsu_single_ecc_error_incr;
	input wire lsu_imprecise_error_load_any;
	input wire lsu_imprecise_error_store_any;
	input wire [31:0] lsu_imprecise_error_addr_any;
	input wire [31:0] exu_div_result;
	input wire exu_div_wren;
	input wire [31:0] exu_csr_rs1_x;
	input wire [31:0] lsu_result_m;
	input wire [31:0] lsu_result_corr_r;
	input wire lsu_load_stall_any;
	input wire lsu_store_stall_any;
	input wire dma_dccm_stall_any;
	input wire dma_iccm_stall_any;
	input wire iccm_dma_sb_error;
	input wire exu_flush_final;
	input wire [31:1] exu_npc_r;
	input wire [31:0] exu_i0_result_x;
	input wire ifu_i0_valid;
	input wire [31:0] ifu_i0_instr;
	input wire [31:1] ifu_i0_pc;
	input wire ifu_i0_pc4;
	input wire [31:1] exu_i0_pc_x;
	input wire mexintpend;
	input wire timer_int;
	input wire soft_int;
	input wire [7:0] pic_claimid;
	input wire [3:0] pic_pl;
	input wire mhwakeup;
	output wire [3:0] dec_tlu_meicurpl;
	output wire [3:0] dec_tlu_meipt;
	input wire [70:0] ifu_ic_debug_rd_data;
	input wire ifu_ic_debug_rd_data_valid;
	output wire [89:0] dec_tlu_ic_diag_pkt;
	input wire dbg_halt_req;
	input wire dbg_resume_req;
	input wire ifu_miss_state_idle;
	output wire dec_tlu_dbg_halted;
	output wire dec_tlu_debug_mode;
	output wire dec_tlu_resume_ack;
	output wire dec_tlu_flush_noredir_r;
	output wire dec_tlu_mpc_halted_only;
	output wire dec_tlu_flush_leak_one_r;
	output wire dec_tlu_flush_err_r;
	output wire [31:2] dec_tlu_meihap;
	output wire dec_debug_wdata_rs1_d;
	output wire [31:0] dec_dbg_rddata;
	output wire dec_dbg_cmd_done;
	output wire dec_dbg_cmd_fail;
	output wire [151:0] trigger_pkt_any;
	output wire dec_tlu_force_halt;
	input wire [1:0] exu_i0_br_hist_r;
	input wire exu_i0_br_error_r;
	input wire exu_i0_br_start_error_r;
	input wire exu_i0_br_valid_r;
	input wire exu_i0_br_mp_r;
	input wire exu_i0_br_middle_r;
	input wire exu_i0_br_way_r;
	output wire dec_i0_rs1_en_d;
	output wire dec_i0_rs2_en_d;
	output wire [31:0] gpr_i0_rs1_d;
	output wire [31:0] gpr_i0_rs2_d;
	output wire [31:0] dec_i0_immed_d;
	output wire [12:1] dec_i0_br_immed_d;
	output wire [43:0] i0_ap;
	output wire dec_i0_alu_decode_d;
	output wire dec_i0_branch_d;
	output wire dec_i0_select_pc_d;
	output wire [31:1] dec_i0_pc_d;
	output wire [3:0] dec_i0_rs1_bypass_en_d;
	output wire [3:0] dec_i0_rs2_bypass_en_d;
	output wire [31:0] dec_i0_result_r;
	output wire [13:0] lsu_p;
	output wire dec_qual_lsu_d;
	output wire [19:0] mul_p;
	output wire [2:0] div_p;
	output wire dec_div_cancel;
	output wire [11:0] dec_lsu_offset_d;
	output wire dec_csr_ren_d;
	output wire [31:0] dec_csr_rddata_d;
	output wire dec_tlu_flush_lower_r;
	output wire dec_tlu_flush_lower_wb;
	output wire [31:1] dec_tlu_flush_path_r;
	output wire dec_tlu_i0_kill_writeb_r;
	output wire dec_tlu_fence_i_r;
	output wire [31:1] pred_correct_npc_x;
	output wire [6:0] dec_tlu_br0_r_pkt;
	output wire dec_tlu_perfcnt0;
	output wire dec_tlu_perfcnt1;
	output wire dec_tlu_perfcnt2;
	output wire dec_tlu_perfcnt3;
	output wire [55:0] dec_i0_predict_p_d;
	output wire [pt[2236-:8] - 1:0] i0_predict_fghr_d;
	output wire [pt[2172-:9]:pt[2163-:6]] i0_predict_index_d;
	output wire [pt[2139-:9] - 1:0] i0_predict_btag_d;
	output wire [$clog2(pt[2061-:14]) - 1:0] dec_fa_error_index;
	output wire dec_lsu_valid_raw_d;
	output wire [31:0] dec_tlu_mrac_ff;
	output wire [1:0] dec_data_en;
	output wire [1:0] dec_ctl_en;
	input wire [15:0] ifu_i0_cinst;
	output wire [103:0] trace_rv_trace_pkt;
	output wire dec_tlu_external_ldfwd_disable;
	output wire dec_tlu_sideeffect_posted_disable;
	output wire dec_tlu_core_ecc_disable;
	output wire dec_tlu_bpred_disable;
	output wire dec_tlu_wb_coalescing_disable;
	output wire [2:0] dec_tlu_dma_qos_prty;
	output wire dec_tlu_misc_clk_override;
	output wire dec_tlu_ifu_clk_override;
	output wire dec_tlu_lsu_clk_override;
	output wire dec_tlu_bus_clk_override;
	output wire dec_tlu_pic_clk_override;
	output wire dec_tlu_picio_clk_override;
	output wire dec_tlu_dccm_clk_override;
	output wire dec_tlu_icm_clk_override;
	output wire dec_tlu_i0_commit_cmt;
	input wire scan_mode;
	wire dec_tlu_dec_clk_override;
	wire clk_override;
	wire dec_ib0_valid_d;
	wire dec_pmu_instr_decoded;
	wire dec_pmu_decode_stall;
	wire dec_pmu_presync_stall;
	wire dec_pmu_postsync_stall;
	wire dec_tlu_wr_pause_r;
	wire [4:0] dec_i0_rs1_d;
	wire [4:0] dec_i0_rs2_d;
	wire [31:0] dec_i0_instr_d;
	wire dec_tlu_trace_disable;
	wire dec_tlu_pipelining_disable;
	wire [4:0] dec_i0_waddr_r;
	wire dec_i0_wen_r;
	wire [31:0] dec_i0_wdata_r;
	wire dec_csr_wen_r;
	wire [11:0] dec_csr_wraddr_r;
	wire [31:0] dec_csr_wrdata_r;
	wire [11:0] dec_csr_rdaddr_d;
	wire dec_csr_legal_d;
	wire dec_csr_wen_unq_d;
	wire dec_csr_any_unq_d;
	wire dec_csr_stall_int_ff;
	wire [16:0] dec_tlu_packet_r;
	wire dec_i0_pc4_d;
	wire dec_tlu_presync_d;
	wire dec_tlu_postsync_d;
	wire dec_tlu_debug_stall;
	wire [31:0] dec_illegal_inst;
	wire dec_i0_icaf_d;
	wire dec_i0_dbecc_d;
	wire dec_i0_icaf_second_d;
	wire [3:0] dec_i0_trigger_match_d;
	wire dec_debug_fence_d;
	wire dec_nonblock_load_wen;
	wire [4:0] dec_nonblock_load_waddr;
	wire dec_tlu_flush_pause_r;
	wire [50:0] dec_i0_brp;
	wire [pt[2172-:9]:pt[2163-:6]] dec_i0_bp_index;
	wire [pt[2236-:8] - 1:0] dec_i0_bp_fghr;
	wire [pt[2139-:9] - 1:0] dec_i0_bp_btag;
	wire [$clog2(pt[2061-:14]) - 1:0] dec_i0_bp_fa_index;
	wire [31:1] dec_tlu_i0_pc_r;
	wire dec_tlu_i0_kill_writeb_wb;
	wire dec_tlu_i0_valid_r;
	wire dec_pause_state;
	wire [1:0] dec_i0_icaf_type_d;
	wire dec_tlu_flush_extint;
	wire [31:0] dec_i0_inst_wb;
	wire [31:1] dec_i0_pc_wb;
	wire dec_tlu_i0_valid_wb1;
	wire dec_tlu_int_valid_wb1;
	wire [4:0] dec_tlu_exc_cause_wb1;
	wire [31:0] dec_tlu_mtval_wb1;
	wire dec_tlu_i0_exc_valid_wb1;
	wire [4:0] div_waddr_wb;
	wire dec_div_active;
	wire dec_debug_valid_d;
	assign clk_override = dec_tlu_dec_clk_override;
	assign dec_dbg_rddata[31:0] = dec_i0_wdata_r[31:0];
	eb1_dec_ib_ctl #(.pt(pt)) instbuff(
		.dbg_cmd_valid(dbg_cmd_valid),
		.dbg_cmd_write(dbg_cmd_write),
		.dbg_cmd_type(dbg_cmd_type),
		.dbg_cmd_addr(dbg_cmd_addr),
		.i0_brp(i0_brp),
		.ifu_i0_bp_index(ifu_i0_bp_index),
		.ifu_i0_bp_fghr(ifu_i0_bp_fghr),
		.ifu_i0_bp_btag(ifu_i0_bp_btag),
		.ifu_i0_fa_index(ifu_i0_fa_index),
		.ifu_i0_pc4(ifu_i0_pc4),
		.ifu_i0_valid(ifu_i0_valid),
		.ifu_i0_icaf(ifu_i0_icaf),
		.ifu_i0_icaf_type(ifu_i0_icaf_type),
		.ifu_i0_icaf_second(ifu_i0_icaf_second),
		.ifu_i0_dbecc(ifu_i0_dbecc),
		.ifu_i0_instr(ifu_i0_instr),
		.ifu_i0_pc(ifu_i0_pc),
		.dec_ib0_valid_d(dec_ib0_valid_d),
		.dec_debug_valid_d(dec_debug_valid_d),
		.dec_i0_instr_d(dec_i0_instr_d),
		.dec_i0_pc_d(dec_i0_pc_d),
		.dec_i0_pc4_d(dec_i0_pc4_d),
		.dec_i0_brp(dec_i0_brp),
		.dec_i0_bp_index(dec_i0_bp_index),
		.dec_i0_bp_fghr(dec_i0_bp_fghr),
		.dec_i0_bp_btag(dec_i0_bp_btag),
		.dec_i0_bp_fa_index(dec_i0_bp_fa_index),
		.dec_i0_icaf_d(dec_i0_icaf_d),
		.dec_i0_icaf_second_d(dec_i0_icaf_second_d),
		.dec_i0_icaf_type_d(dec_i0_icaf_type_d),
		.dec_i0_dbecc_d(dec_i0_dbecc_d),
		.dec_debug_wdata_rs1_d(dec_debug_wdata_rs1_d),
		.dec_debug_fence_d(dec_debug_fence_d)
	);
	eb1_dec_decode_ctl #(.pt(pt)) decode(
		.dec_tlu_trace_disable(dec_tlu_trace_disable),
		.dec_debug_valid_d(dec_debug_valid_d),
		.dec_tlu_flush_extint(dec_tlu_flush_extint),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.dec_extint_stall(dec_extint_stall),
		.ifu_i0_cinst(ifu_i0_cinst),
		.dec_i0_inst_wb(dec_i0_inst_wb),
		.dec_i0_pc_wb(dec_i0_pc_wb),
		.lsu_nonblock_load_valid_m(lsu_nonblock_load_valid_m),
		.lsu_nonblock_load_tag_m(lsu_nonblock_load_tag_m),
		.lsu_nonblock_load_inv_r(lsu_nonblock_load_inv_r),
		.lsu_nonblock_load_inv_tag_r(lsu_nonblock_load_inv_tag_r),
		.lsu_nonblock_load_data_valid(lsu_nonblock_load_data_valid),
		.lsu_nonblock_load_data_error(lsu_nonblock_load_data_error),
		.lsu_nonblock_load_data_tag(lsu_nonblock_load_data_tag),
		.dec_i0_trigger_match_d(dec_i0_trigger_match_d),
		.dec_tlu_wr_pause_r(dec_tlu_wr_pause_r),
		.dec_tlu_pipelining_disable(dec_tlu_pipelining_disable),
		.lsu_trigger_match_m(lsu_trigger_match_m),
		.lsu_pmu_misaligned_m(lsu_pmu_misaligned_m),
		.dec_tlu_debug_stall(dec_tlu_debug_stall),
		.dec_tlu_flush_leak_one_r(dec_tlu_flush_leak_one_r),
		.dec_debug_fence_d(dec_debug_fence_d),
		.dbg_cmd_wrdata(dbg_cmd_wrdata),
		.dec_i0_icaf_d(dec_i0_icaf_d),
		.dec_i0_icaf_second_d(dec_i0_icaf_second_d),
		.dec_i0_icaf_type_d(dec_i0_icaf_type_d),
		.dec_i0_dbecc_d(dec_i0_dbecc_d),
		.dec_i0_brp(dec_i0_brp),
		.dec_i0_bp_index(dec_i0_bp_index),
		.dec_i0_bp_fghr(dec_i0_bp_fghr),
		.dec_i0_bp_btag(dec_i0_bp_btag),
		.dec_i0_bp_fa_index(dec_i0_bp_fa_index),
		.lsu_idle_any(lsu_idle_any),
		.lsu_load_stall_any(lsu_load_stall_any),
		.lsu_store_stall_any(lsu_store_stall_any),
		.dma_dccm_stall_any(dma_dccm_stall_any),
		.exu_div_wren(exu_div_wren),
		.dec_tlu_i0_kill_writeb_wb(dec_tlu_i0_kill_writeb_wb),
		.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_wb),
		.dec_tlu_i0_kill_writeb_r(dec_tlu_i0_kill_writeb_r),
		.dec_tlu_flush_lower_r(dec_tlu_flush_lower_r),
		.dec_tlu_flush_pause_r(dec_tlu_flush_pause_r),
		.dec_tlu_presync_d(dec_tlu_presync_d),
		.dec_tlu_postsync_d(dec_tlu_postsync_d),
		.dec_i0_pc4_d(dec_i0_pc4_d),
		.dec_csr_rddata_d(dec_csr_rddata_d),
		.dec_csr_legal_d(dec_csr_legal_d),
		.exu_csr_rs1_x(exu_csr_rs1_x),
		.lsu_result_m(lsu_result_m),
		.lsu_result_corr_r(lsu_result_corr_r),
		.exu_flush_final(exu_flush_final),
		.exu_i0_pc_x(exu_i0_pc_x),
		.dec_i0_instr_d(dec_i0_instr_d),
		.dec_ib0_valid_d(dec_ib0_valid_d),
		.exu_i0_result_x(exu_i0_result_x),
		.clk(clk),
		.active_clk(active_clk),
		.free_l2clk(free_l2clk),
		.clk_override(clk_override),
		.rst_l(rst_l),
		.dec_i0_rs1_en_d(dec_i0_rs1_en_d),
		.dec_i0_rs2_en_d(dec_i0_rs2_en_d),
		.dec_i0_rs1_d(dec_i0_rs1_d),
		.dec_i0_rs2_d(dec_i0_rs2_d),
		.dec_i0_immed_d(dec_i0_immed_d),
		.dec_i0_br_immed_d(dec_i0_br_immed_d),
		.i0_ap(i0_ap),
		.dec_i0_decode_d(dec_i0_decode_d),
		.dec_i0_alu_decode_d(dec_i0_alu_decode_d),
		.dec_i0_branch_d(dec_i0_branch_d),
		.dec_i0_waddr_r(dec_i0_waddr_r),
		.dec_i0_wen_r(dec_i0_wen_r),
		.dec_i0_wdata_r(dec_i0_wdata_r),
		.dec_i0_select_pc_d(dec_i0_select_pc_d),
		.dec_i0_rs1_bypass_en_d(dec_i0_rs1_bypass_en_d),
		.dec_i0_rs2_bypass_en_d(dec_i0_rs2_bypass_en_d),
		.dec_i0_result_r(dec_i0_result_r),
		.lsu_p(lsu_p),
		.dec_qual_lsu_d(dec_qual_lsu_d),
		.mul_p(mul_p),
		.div_p(div_p),
		.div_waddr_wb(div_waddr_wb),
		.dec_div_cancel(dec_div_cancel),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.dec_lsu_offset_d(dec_lsu_offset_d),
		.dec_csr_ren_d(dec_csr_ren_d),
		.dec_csr_wen_unq_d(dec_csr_wen_unq_d),
		.dec_csr_any_unq_d(dec_csr_any_unq_d),
		.dec_csr_rdaddr_d(dec_csr_rdaddr_d),
		.dec_csr_wen_r(dec_csr_wen_r),
		.dec_csr_wraddr_r(dec_csr_wraddr_r),
		.dec_csr_wrdata_r(dec_csr_wrdata_r),
		.dec_csr_stall_int_ff(dec_csr_stall_int_ff),
		.dec_tlu_i0_valid_r(dec_tlu_i0_valid_r),
		.dec_tlu_packet_r(dec_tlu_packet_r),
		.dec_tlu_i0_pc_r(dec_tlu_i0_pc_r),
		.dec_illegal_inst(dec_illegal_inst),
		.pred_correct_npc_x(pred_correct_npc_x),
		.dec_i0_predict_p_d(dec_i0_predict_p_d),
		.i0_predict_fghr_d(i0_predict_fghr_d),
		.i0_predict_index_d(i0_predict_index_d),
		.i0_predict_btag_d(i0_predict_btag_d),
		.dec_fa_error_index(dec_fa_error_index),
		.dec_data_en(dec_data_en),
		.dec_ctl_en(dec_ctl_en),
		.dec_pmu_instr_decoded(dec_pmu_instr_decoded),
		.dec_pmu_decode_stall(dec_pmu_decode_stall),
		.dec_pmu_presync_stall(dec_pmu_presync_stall),
		.dec_pmu_postsync_stall(dec_pmu_postsync_stall),
		.dec_nonblock_load_wen(dec_nonblock_load_wen),
		.dec_nonblock_load_waddr(dec_nonblock_load_waddr),
		.dec_pause_state(dec_pause_state),
		.dec_pause_state_cg(dec_pause_state_cg),
		.dec_div_active(dec_div_active),
		.scan_mode(scan_mode)
	);
	eb1_dec_tlu_ctl #(.pt(pt)) tlu(
		.clk(clk),
		.free_clk(free_clk),
		.free_l2clk(free_l2clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.rst_vec(rst_vec),
		.nmi_int(nmi_int),
		.nmi_vec(nmi_vec),
		.i_cpu_halt_req(i_cpu_halt_req),
		.i_cpu_run_req(i_cpu_run_req),
		.lsu_fastint_stall_any(lsu_fastint_stall_any),
		.ifu_pmu_instr_aligned(ifu_pmu_instr_aligned),
		.ifu_pmu_fetch_stall(ifu_pmu_fetch_stall),
		.ifu_pmu_ic_miss(ifu_pmu_ic_miss),
		.ifu_pmu_ic_hit(ifu_pmu_ic_hit),
		.ifu_pmu_bus_error(ifu_pmu_bus_error),
		.ifu_pmu_bus_busy(ifu_pmu_bus_busy),
		.ifu_pmu_bus_trxn(ifu_pmu_bus_trxn),
		.dec_pmu_instr_decoded(dec_pmu_instr_decoded),
		.dec_pmu_decode_stall(dec_pmu_decode_stall),
		.dec_pmu_presync_stall(dec_pmu_presync_stall),
		.dec_pmu_postsync_stall(dec_pmu_postsync_stall),
		.lsu_store_stall_any(lsu_store_stall_any),
		.dma_dccm_stall_any(dma_dccm_stall_any),
		.dma_iccm_stall_any(dma_iccm_stall_any),
		.exu_pmu_i0_br_misp(exu_pmu_i0_br_misp),
		.exu_pmu_i0_br_ataken(exu_pmu_i0_br_ataken),
		.exu_pmu_i0_pc4(exu_pmu_i0_pc4),
		.lsu_pmu_bus_trxn(lsu_pmu_bus_trxn),
		.lsu_pmu_bus_misaligned(lsu_pmu_bus_misaligned),
		.lsu_pmu_bus_error(lsu_pmu_bus_error),
		.lsu_pmu_bus_busy(lsu_pmu_bus_busy),
		.lsu_pmu_load_external_m(lsu_pmu_load_external_m),
		.lsu_pmu_store_external_m(lsu_pmu_store_external_m),
		.dma_pmu_dccm_read(dma_pmu_dccm_read),
		.dma_pmu_dccm_write(dma_pmu_dccm_write),
		.dma_pmu_any_read(dma_pmu_any_read),
		.dma_pmu_any_write(dma_pmu_any_write),
		.lsu_fir_addr(lsu_fir_addr),
		.lsu_fir_error(lsu_fir_error),
		.iccm_dma_sb_error(iccm_dma_sb_error),
		.lsu_error_pkt_r(lsu_error_pkt_r),
		.lsu_single_ecc_error_incr(lsu_single_ecc_error_incr),
		.dec_pause_state(dec_pause_state),
		.lsu_imprecise_error_store_any(lsu_imprecise_error_store_any),
		.lsu_imprecise_error_load_any(lsu_imprecise_error_load_any),
		.lsu_imprecise_error_addr_any(lsu_imprecise_error_addr_any),
		.dec_csr_wen_unq_d(dec_csr_wen_unq_d),
		.dec_csr_any_unq_d(dec_csr_any_unq_d),
		.dec_csr_rdaddr_d(dec_csr_rdaddr_d),
		.dec_csr_wen_r(dec_csr_wen_r),
		.dec_csr_wraddr_r(dec_csr_wraddr_r),
		.dec_csr_wrdata_r(dec_csr_wrdata_r),
		.dec_csr_stall_int_ff(dec_csr_stall_int_ff),
		.dec_tlu_i0_valid_r(dec_tlu_i0_valid_r),
		.exu_npc_r(exu_npc_r),
		.dec_tlu_i0_pc_r(dec_tlu_i0_pc_r),
		.dec_tlu_packet_r(dec_tlu_packet_r),
		.dec_illegal_inst(dec_illegal_inst),
		.dec_i0_decode_d(dec_i0_decode_d),
		.exu_i0_br_hist_r(exu_i0_br_hist_r),
		.exu_i0_br_error_r(exu_i0_br_error_r),
		.exu_i0_br_start_error_r(exu_i0_br_start_error_r),
		.exu_i0_br_valid_r(exu_i0_br_valid_r),
		.exu_i0_br_mp_r(exu_i0_br_mp_r),
		.exu_i0_br_middle_r(exu_i0_br_middle_r),
		.exu_i0_br_way_r(exu_i0_br_way_r),
		.dec_tlu_core_empty(dec_tlu_core_empty),
		.dec_dbg_cmd_done(dec_dbg_cmd_done),
		.dec_dbg_cmd_fail(dec_dbg_cmd_fail),
		.dec_tlu_dbg_halted(dec_tlu_dbg_halted),
		.dec_tlu_debug_mode(dec_tlu_debug_mode),
		.dec_tlu_resume_ack(dec_tlu_resume_ack),
		.dec_tlu_debug_stall(dec_tlu_debug_stall),
		.dec_tlu_flush_noredir_r(dec_tlu_flush_noredir_r),
		.dec_tlu_mpc_halted_only(dec_tlu_mpc_halted_only),
		.dec_tlu_flush_leak_one_r(dec_tlu_flush_leak_one_r),
		.dec_tlu_flush_err_r(dec_tlu_flush_err_r),
		.dec_tlu_flush_extint(dec_tlu_flush_extint),
		.dec_tlu_meihap(dec_tlu_meihap),
		.dbg_halt_req(dbg_halt_req),
		.dbg_resume_req(dbg_resume_req),
		.ifu_miss_state_idle(ifu_miss_state_idle),
		.lsu_idle_any(lsu_idle_any),
		.dec_div_active(dec_div_active),
		.trigger_pkt_any(trigger_pkt_any),
		.ifu_ic_error_start(ifu_ic_error_start),
		.ifu_iccm_rd_ecc_single_err(ifu_iccm_rd_ecc_single_err),
		.ifu_ic_debug_rd_data(ifu_ic_debug_rd_data),
		.ifu_ic_debug_rd_data_valid(ifu_ic_debug_rd_data_valid),
		.dec_tlu_ic_diag_pkt(dec_tlu_ic_diag_pkt),
		.pic_claimid(pic_claimid),
		.pic_pl(pic_pl),
		.mhwakeup(mhwakeup),
		.mexintpend(mexintpend),
		.timer_int(timer_int),
		.soft_int(soft_int),
		.o_cpu_halt_status(o_cpu_halt_status),
		.o_cpu_halt_ack(o_cpu_halt_ack),
		.o_cpu_run_ack(o_cpu_run_ack),
		.o_debug_mode_status(o_debug_mode_status),
		.core_id(core_id),
		.mpc_debug_halt_req(mpc_debug_halt_req),
		.mpc_debug_run_req(mpc_debug_run_req),
		.mpc_reset_run_req(mpc_reset_run_req),
		.mpc_debug_halt_ack(mpc_debug_halt_ack),
		.mpc_debug_run_ack(mpc_debug_run_ack),
		.debug_brkpt_status(debug_brkpt_status),
		.dec_tlu_meicurpl(dec_tlu_meicurpl),
		.dec_tlu_meipt(dec_tlu_meipt),
		.dec_csr_rddata_d(dec_csr_rddata_d),
		.dec_csr_legal_d(dec_csr_legal_d),
		.dec_tlu_br0_r_pkt(dec_tlu_br0_r_pkt),
		.dec_tlu_i0_kill_writeb_wb(dec_tlu_i0_kill_writeb_wb),
		.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_wb),
		.dec_tlu_i0_commit_cmt(dec_tlu_i0_commit_cmt),
		.dec_tlu_i0_kill_writeb_r(dec_tlu_i0_kill_writeb_r),
		.dec_tlu_flush_lower_r(dec_tlu_flush_lower_r),
		.dec_tlu_flush_path_r(dec_tlu_flush_path_r),
		.dec_tlu_fence_i_r(dec_tlu_fence_i_r),
		.dec_tlu_wr_pause_r(dec_tlu_wr_pause_r),
		.dec_tlu_flush_pause_r(dec_tlu_flush_pause_r),
		.dec_tlu_presync_d(dec_tlu_presync_d),
		.dec_tlu_postsync_d(dec_tlu_postsync_d),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.dec_tlu_perfcnt0(dec_tlu_perfcnt0),
		.dec_tlu_perfcnt1(dec_tlu_perfcnt1),
		.dec_tlu_perfcnt2(dec_tlu_perfcnt2),
		.dec_tlu_perfcnt3(dec_tlu_perfcnt3),
		.dec_tlu_i0_exc_valid_wb1(dec_tlu_i0_exc_valid_wb1),
		.dec_tlu_i0_valid_wb1(dec_tlu_i0_valid_wb1),
		.dec_tlu_int_valid_wb1(dec_tlu_int_valid_wb1),
		.dec_tlu_exc_cause_wb1(dec_tlu_exc_cause_wb1),
		.dec_tlu_mtval_wb1(dec_tlu_mtval_wb1),
		.dec_tlu_external_ldfwd_disable(dec_tlu_external_ldfwd_disable),
		.dec_tlu_sideeffect_posted_disable(dec_tlu_sideeffect_posted_disable),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.dec_tlu_bpred_disable(dec_tlu_bpred_disable),
		.dec_tlu_wb_coalescing_disable(dec_tlu_wb_coalescing_disable),
		.dec_tlu_pipelining_disable(dec_tlu_pipelining_disable),
		.dec_tlu_trace_disable(dec_tlu_trace_disable),
		.dec_tlu_dma_qos_prty(dec_tlu_dma_qos_prty),
		.dec_tlu_misc_clk_override(dec_tlu_misc_clk_override),
		.dec_tlu_dec_clk_override(dec_tlu_dec_clk_override),
		.dec_tlu_ifu_clk_override(dec_tlu_ifu_clk_override),
		.dec_tlu_lsu_clk_override(dec_tlu_lsu_clk_override),
		.dec_tlu_bus_clk_override(dec_tlu_bus_clk_override),
		.dec_tlu_pic_clk_override(dec_tlu_pic_clk_override),
		.dec_tlu_picio_clk_override(dec_tlu_picio_clk_override),
		.dec_tlu_dccm_clk_override(dec_tlu_dccm_clk_override),
		.dec_tlu_icm_clk_override(dec_tlu_icm_clk_override)
	);
	eb1_dec_gpr_ctl #(.pt(pt)) arf(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.raddr0(dec_i0_rs1_d[4:0]),
		.raddr1(dec_i0_rs2_d[4:0]),
		.wen0(dec_i0_wen_r),
		.waddr0(dec_i0_waddr_r[4:0]),
		.wd0(dec_i0_wdata_r[31:0]),
		.wen1(dec_nonblock_load_wen),
		.waddr1(dec_nonblock_load_waddr[4:0]),
		.wd1(lsu_nonblock_load_data[31:0]),
		.wen2(exu_div_wren),
		.waddr2(div_waddr_wb),
		.wd2(exu_div_result[31:0]),
		.rd0(gpr_i0_rs1_d[31:0]),
		.rd1(gpr_i0_rs2_d[31:0])
	);
	eb1_dec_trigger #(.pt(pt)) dec_trigger(
		.trigger_pkt_any(trigger_pkt_any),
		.dec_i0_pc_d(dec_i0_pc_d),
		.dec_i0_trigger_match_d(dec_i0_trigger_match_d)
	);
	assign trace_rv_trace_pkt[102-:32] = dec_i0_inst_wb[31:0];
	assign trace_rv_trace_pkt[70-:32] = {dec_i0_pc_wb[31:1], 1'b0};
	assign trace_rv_trace_pkt[103] = (dec_tlu_int_valid_wb1 | dec_tlu_i0_valid_wb1) | dec_tlu_i0_exc_valid_wb1;
	assign trace_rv_trace_pkt[38] = dec_tlu_int_valid_wb1 | dec_tlu_i0_exc_valid_wb1;
	assign trace_rv_trace_pkt[37-:5] = dec_tlu_exc_cause_wb1[4:0];
	assign trace_rv_trace_pkt[32] = dec_tlu_int_valid_wb1;
	assign trace_rv_trace_pkt[31-:32] = dec_tlu_mtval_wb1[31:0];
endmodule
module eb1_dec_decode_ctl (
	dec_tlu_trace_disable,
	dec_debug_valid_d,
	dec_tlu_flush_extint,
	dec_tlu_force_halt,
	dec_extint_stall,
	ifu_i0_cinst,
	dec_i0_inst_wb,
	dec_i0_pc_wb,
	lsu_nonblock_load_valid_m,
	lsu_nonblock_load_tag_m,
	lsu_nonblock_load_inv_r,
	lsu_nonblock_load_inv_tag_r,
	lsu_nonblock_load_data_valid,
	lsu_nonblock_load_data_error,
	lsu_nonblock_load_data_tag,
	dec_i0_trigger_match_d,
	dec_tlu_wr_pause_r,
	dec_tlu_pipelining_disable,
	lsu_trigger_match_m,
	lsu_pmu_misaligned_m,
	dec_tlu_debug_stall,
	dec_tlu_flush_leak_one_r,
	dec_debug_fence_d,
	dbg_cmd_wrdata,
	dec_i0_icaf_d,
	dec_i0_icaf_second_d,
	dec_i0_icaf_type_d,
	dec_i0_dbecc_d,
	dec_i0_brp,
	dec_i0_bp_index,
	dec_i0_bp_fghr,
	dec_i0_bp_btag,
	dec_i0_bp_fa_index,
	lsu_idle_any,
	lsu_load_stall_any,
	lsu_store_stall_any,
	dma_dccm_stall_any,
	exu_div_wren,
	dec_tlu_i0_kill_writeb_wb,
	dec_tlu_flush_lower_wb,
	dec_tlu_i0_kill_writeb_r,
	dec_tlu_flush_lower_r,
	dec_tlu_flush_pause_r,
	dec_tlu_presync_d,
	dec_tlu_postsync_d,
	dec_i0_pc4_d,
	dec_csr_rddata_d,
	dec_csr_legal_d,
	exu_csr_rs1_x,
	lsu_result_m,
	lsu_result_corr_r,
	exu_flush_final,
	exu_i0_pc_x,
	dec_i0_instr_d,
	dec_ib0_valid_d,
	exu_i0_result_x,
	clk,
	active_clk,
	free_l2clk,
	clk_override,
	rst_l,
	dec_i0_rs1_en_d,
	dec_i0_rs2_en_d,
	dec_i0_rs1_d,
	dec_i0_rs2_d,
	dec_i0_immed_d,
	dec_i0_br_immed_d,
	i0_ap,
	dec_i0_decode_d,
	dec_i0_alu_decode_d,
	dec_i0_branch_d,
	dec_i0_waddr_r,
	dec_i0_wen_r,
	dec_i0_wdata_r,
	dec_i0_select_pc_d,
	dec_i0_rs1_bypass_en_d,
	dec_i0_rs2_bypass_en_d,
	dec_i0_result_r,
	lsu_p,
	dec_qual_lsu_d,
	mul_p,
	div_p,
	div_waddr_wb,
	dec_div_cancel,
	dec_lsu_valid_raw_d,
	dec_lsu_offset_d,
	dec_csr_ren_d,
	dec_csr_wen_unq_d,
	dec_csr_any_unq_d,
	dec_csr_rdaddr_d,
	dec_csr_wen_r,
	dec_csr_wraddr_r,
	dec_csr_wrdata_r,
	dec_csr_stall_int_ff,
	dec_tlu_i0_valid_r,
	dec_tlu_packet_r,
	dec_tlu_i0_pc_r,
	dec_illegal_inst,
	pred_correct_npc_x,
	dec_i0_predict_p_d,
	i0_predict_fghr_d,
	i0_predict_index_d,
	i0_predict_btag_d,
	dec_fa_error_index,
	dec_data_en,
	dec_ctl_en,
	dec_pmu_instr_decoded,
	dec_pmu_decode_stall,
	dec_pmu_presync_stall,
	dec_pmu_postsync_stall,
	dec_nonblock_load_wen,
	dec_nonblock_load_waddr,
	dec_pause_state,
	dec_pause_state_cg,
	dec_div_active,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire dec_tlu_trace_disable;
	input wire dec_debug_valid_d;
	input wire dec_tlu_flush_extint;
	input wire dec_tlu_force_halt;
	output wire dec_extint_stall;
	input wire [15:0] ifu_i0_cinst;
	output wire [31:0] dec_i0_inst_wb;
	output wire [31:1] dec_i0_pc_wb;
	input wire lsu_nonblock_load_valid_m;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	input wire lsu_nonblock_load_inv_r;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	input wire lsu_nonblock_load_data_valid;
	input wire lsu_nonblock_load_data_error;
	input wire [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	input wire [3:0] dec_i0_trigger_match_d;
	input wire dec_tlu_wr_pause_r;
	input wire dec_tlu_pipelining_disable;
	input wire [3:0] lsu_trigger_match_m;
	input wire lsu_pmu_misaligned_m;
	input wire dec_tlu_debug_stall;
	input wire dec_tlu_flush_leak_one_r;
	input wire dec_debug_fence_d;
	input wire [1:0] dbg_cmd_wrdata;
	input wire dec_i0_icaf_d;
	input wire dec_i0_icaf_second_d;
	input wire [1:0] dec_i0_icaf_type_d;
	input wire dec_i0_dbecc_d;
	input wire [50:0] dec_i0_brp;
	input wire [pt[2172-:9]:pt[2163-:6]] dec_i0_bp_index;
	input wire [pt[2236-:8] - 1:0] dec_i0_bp_fghr;
	input wire [pt[2139-:9] - 1:0] dec_i0_bp_btag;
	input wire [$clog2(pt[2061-:14]) - 1:0] dec_i0_bp_fa_index;
	input wire lsu_idle_any;
	input wire lsu_load_stall_any;
	input wire lsu_store_stall_any;
	input wire dma_dccm_stall_any;
	input wire exu_div_wren;
	input wire dec_tlu_i0_kill_writeb_wb;
	input wire dec_tlu_flush_lower_wb;
	input wire dec_tlu_i0_kill_writeb_r;
	input wire dec_tlu_flush_lower_r;
	input wire dec_tlu_flush_pause_r;
	input wire dec_tlu_presync_d;
	input wire dec_tlu_postsync_d;
	input wire dec_i0_pc4_d;
	input wire [31:0] dec_csr_rddata_d;
	input wire dec_csr_legal_d;
	input wire [31:0] exu_csr_rs1_x;
	input wire [31:0] lsu_result_m;
	input wire [31:0] lsu_result_corr_r;
	input wire exu_flush_final;
	input wire [31:1] exu_i0_pc_x;
	input wire [31:0] dec_i0_instr_d;
	input wire dec_ib0_valid_d;
	input wire [31:0] exu_i0_result_x;
	input wire clk;
	input wire active_clk;
	input wire free_l2clk;
	input wire clk_override;
	input wire rst_l;
	output wire dec_i0_rs1_en_d;
	output wire dec_i0_rs2_en_d;
	output wire [4:0] dec_i0_rs1_d;
	output wire [4:0] dec_i0_rs2_d;
	output wire [31:0] dec_i0_immed_d;
	output wire [12:1] dec_i0_br_immed_d;
	output wire [43:0] i0_ap;
	output wire dec_i0_decode_d;
	output wire dec_i0_alu_decode_d;
	output wire dec_i0_branch_d;
	output wire [4:0] dec_i0_waddr_r;
	output wire dec_i0_wen_r;
	output wire [31:0] dec_i0_wdata_r;
	output wire dec_i0_select_pc_d;
	output wire [3:0] dec_i0_rs1_bypass_en_d;
	output wire [3:0] dec_i0_rs2_bypass_en_d;
	output wire [31:0] dec_i0_result_r;
	output reg [13:0] lsu_p;
	output wire dec_qual_lsu_d;
	output wire [19:0] mul_p;
	output wire [2:0] div_p;
	output wire [4:0] div_waddr_wb;
	output wire dec_div_cancel;
	output wire dec_lsu_valid_raw_d;
	output wire [11:0] dec_lsu_offset_d;
	output wire dec_csr_ren_d;
	output wire dec_csr_wen_unq_d;
	output wire dec_csr_any_unq_d;
	output wire [11:0] dec_csr_rdaddr_d;
	output wire dec_csr_wen_r;
	output wire [11:0] dec_csr_wraddr_r;
	output wire [31:0] dec_csr_wrdata_r;
	output wire dec_csr_stall_int_ff;
	output dec_tlu_i0_valid_r;
	output reg [16:0] dec_tlu_packet_r;
	output wire [31:1] dec_tlu_i0_pc_r;
	output wire [31:0] dec_illegal_inst;
	output wire [31:1] pred_correct_npc_x;
	output reg [55:0] dec_i0_predict_p_d;
	output wire [pt[2236-:8] - 1:0] i0_predict_fghr_d;
	output wire [pt[2172-:9]:pt[2163-:6]] i0_predict_index_d;
	output wire [pt[2139-:9] - 1:0] i0_predict_btag_d;
	output wire [$clog2(pt[2061-:14]) - 1:0] dec_fa_error_index;
	output wire [1:0] dec_data_en;
	output wire [1:0] dec_ctl_en;
	output wire dec_pmu_instr_decoded;
	output wire dec_pmu_decode_stall;
	output wire dec_pmu_presync_stall;
	output wire dec_pmu_postsync_stall;
	output wire dec_nonblock_load_wen;
	output reg [4:0] dec_nonblock_load_waddr;
	output wire dec_pause_state;
	output wire dec_pause_state_cg;
	output wire dec_div_active;
	input wire scan_mode;
	wire [94:0] i0_dp_raw;
	reg [94:0] i0_dp;
	wire [31:0] i0;
	wire i0_valid_d;
	wire [31:0] i0_result_r;
	wire [2:0] i0_rs1bypass;
	wire [2:0] i0_rs2bypass;
	wire i0_jalimm20;
	wire i0_uiimm20;
	wire lsu_decode_d;
	wire [31:0] i0_immed_d;
	wire i0_presync;
	wire i0_postsync;
	wire postsync_stall;
	wire ps_stall;
	wire prior_inflight;
	wire prior_inflight_wb;
	wire csr_clr_d;
	wire csr_set_d;
	wire csr_write_d;
	wire csr_clr_x;
	wire csr_set_x;
	wire csr_write_x;
	wire csr_imm_x;
	wire [31:0] csr_mask_x;
	wire [31:0] write_csr_data_x;
	wire [31:0] write_csr_data_in;
	wire [31:0] write_csr_data;
	wire csr_data_wen;
	wire [4:0] csrimm_x;
	wire [31:0] csr_rddata_x;
	wire mul_decode_d;
	wire div_decode_d;
	wire div_e1_to_r;
	wire div_flush;
	wire div_active_in;
	wire div_active;
	wire i0_nonblock_div_stall;
	wire i0_div_prior_div_stall;
	wire nonblock_div_cancel;
	wire i0_legal;
	wire shift_illegal;
	wire illegal_inst_en;
	wire illegal_lockout_in;
	wire illegal_lockout;
	wire i0_legal_decode_d;
	wire i0_exulegal_decode_d;
	wire i0_exudecode_d;
	wire i0_exublock_d;
	wire [12:1] last_br_immed_d;
	wire i0_rs1_depend_i0_x;
	wire i0_rs1_depend_i0_r;
	wire i0_rs2_depend_i0_x;
	wire i0_rs2_depend_i0_r;
	wire i0_div_decode_d;
	wire i0_load_block_d;
	wire [1:0] i0_rs1_depth_d;
	wire [1:0] i0_rs2_depth_d;
	wire i0_load_stall_d;
	wire i0_store_stall_d;
	wire i0_predict_nt;
	wire i0_predict_t;
	wire i0_notbr_error;
	wire i0_br_toffset_error;
	wire i0_ret_error;
	wire i0_br_error;
	wire i0_br_error_all;
	wire [11:0] i0_br_offset;
	wire [20:1] i0_pcall_imm;
	wire i0_pcall_12b_offset;
	wire i0_pcall_raw;
	wire i0_pcall_case;
	wire i0_pcall;
	wire i0_pja_raw;
	wire i0_pja_case;
	wire i0_pja;
	wire i0_pret_case;
	wire i0_pret_raw;
	wire i0_pret;
	wire i0_jal;
	wire i0_predict_br;
	wire store_data_bypass_d;
	wire store_data_bypass_m;
	wire [2:0] i0_rs1_class_d;
	wire [2:0] i0_rs2_class_d;
	wire [2:0] i0_d_c;
	wire [2:0] i0_x_c;
	wire [2:0] i0_r_c;
	wire i0_ap_pc2;
	wire i0_ap_pc4;
	wire i0_rd_en_d;
	wire load_ldst_bypass_d;
	wire leak1_i0_stall_in;
	wire leak1_i0_stall;
	wire leak1_i1_stall_in;
	wire leak1_i1_stall;
	wire leak1_mode;
	wire i0_csr_write_only_d;
	wire prior_inflight_x;
	wire prior_inflight_eff;
	wire any_csr_d;
	wire prior_csr_write;
	wire [3:0] i0_pipe_en;
	wire i0_r_ctl_en;
	wire i0_x_ctl_en;
	wire i0_wb_ctl_en;
	wire i0_x_data_en;
	wire i0_r_data_en;
	wire i0_wb_data_en;
	wire debug_fence_i;
	wire debug_fence;
	wire i0_csr_write;
	wire presync_stall;
	wire i0_instr_error;
	wire i0_icaf_d;
	wire clear_pause;
	wire pause_state_in;
	wire pause_state;
	wire pause_stall;
	wire i0_brp_valid;
	wire nonblock_load_cancel;
	wire lsu_idle;
	wire lsu_pmu_misaligned_r;
	wire csr_ren_qual_d;
	wire csr_read_x;
	wire i0_block_d;
	wire i0_block_raw_d;
	wire ps_stall_in;
	wire [31:0] i0_result_x;
	wire [23:0] d_d;
	wire [23:0] x_d;
	wire [23:0] r_d;
	wire [23:0] wbd;
	reg [23:0] x_d_in;
	reg [23:0] r_d_in;
	wire [16:0] d_t;
	wire [16:0] x_t;
	reg [16:0] x_t_in;
	reg [16:0] r_t_in;
	wire [16:0] r_t;
	wire [3:0] lsu_trigger_match_r;
	wire [31:1] dec_i0_pc_r;
	wire csr_read;
	wire csr_write;
	wire i0_br_unpred;
	wire nonblock_load_valid_m_delay;
	wire i0_wen_r;
	wire tlu_wr_pause_r1;
	wire tlu_wr_pause_r2;
	wire flush_final_r;
	wire bitmanip_zbb_legal;
	wire bitmanip_zbs_legal;
	wire bitmanip_zbe_legal;
	wire bitmanip_zbc_legal;
	wire bitmanip_zbp_legal;
	wire bitmanip_zbr_legal;
	wire bitmanip_zbf_legal;
	wire bitmanip_zba_legal;
	wire bitmanip_zbb_zbp_legal;
	wire bitmanip_legal;
	wire data_gate_en;
	wire data_gate_clk;
	localparam NBLOAD_SIZE = pt[173-:9];
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	localparam NBLOAD_SIZE_MSB = sv2v_cast_32_signed(pt[173-:9]) - 1;
	localparam NBLOAD_TAG_MSB = pt[164-:7] - 1;
	wire cam_write;
	wire cam_inv_reset;
	wire cam_data_reset;
	wire [NBLOAD_TAG_MSB:0] cam_write_tag;
	wire [NBLOAD_TAG_MSB:0] cam_inv_reset_tag;
	wire [NBLOAD_TAG_MSB:0] cam_data_reset_tag;
	reg [NBLOAD_SIZE_MSB:0] cam_wen;
	wire [NBLOAD_TAG_MSB:0] load_data_tag;
	wire [NBLOAD_SIZE_MSB:0] nonblock_load_write;
	reg [(NBLOAD_SIZE_MSB >= 0 ? ((NBLOAD_SIZE_MSB + 1) * 10) - 1 : ((1 - NBLOAD_SIZE_MSB) * 10) + ((NBLOAD_SIZE_MSB * 10) - 1)):(NBLOAD_SIZE_MSB >= 0 ? 0 : NBLOAD_SIZE_MSB * 10)] cam;
	reg [(NBLOAD_SIZE_MSB >= 0 ? ((NBLOAD_SIZE_MSB + 1) * 10) - 1 : ((1 - NBLOAD_SIZE_MSB) * 10) + ((NBLOAD_SIZE_MSB * 10) - 1)):(NBLOAD_SIZE_MSB >= 0 ? 0 : NBLOAD_SIZE_MSB * 10)] cam_in;
	wire [(NBLOAD_SIZE_MSB >= 0 ? ((NBLOAD_SIZE_MSB + 1) * 10) - 1 : ((1 - NBLOAD_SIZE_MSB) * 10) + ((NBLOAD_SIZE_MSB * 10) - 1)):(NBLOAD_SIZE_MSB >= 0 ? 0 : NBLOAD_SIZE_MSB * 10)] cam_raw;
	wire [4:0] nonblock_load_rd;
	reg i0_nonblock_load_stall;
	wire i0_nonblock_boundary_stall;
	wire i0_rs1_nonblock_load_bypass_en_d;
	wire i0_rs2_nonblock_load_bypass_en_d;
	wire i0_load_kill_wen_r;
	reg found;
	wire [NBLOAD_SIZE_MSB:0] cam_inv_reset_val;
	wire [NBLOAD_SIZE_MSB:0] cam_data_reset_val;
	wire debug_fence_raw;
	wire [31:0] i0_result_r_raw;
	wire [31:0] i0_result_corr_r;
	wire [12:1] last_br_immed_x;
	wire [31:0] i0_inst_d;
	wire [31:0] i0_inst_x;
	wire [31:0] i0_inst_r;
	wire [31:0] i0_inst_wb_in;
	wire [31:0] i0_inst_wb;
	wire [31:1] i0_pc_wb;
	wire i0_wb_en;
	wire trace_enable;
	wire debug_valid_x;
	reg [3:0] i0_itype;
	wire [14:0] i0r;
	rvdffie #(.WIDTH(8)) misc1ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({leak1_i1_stall_in, leak1_i0_stall_in, dec_tlu_flush_extint, pause_state_in, dec_tlu_wr_pause_r, tlu_wr_pause_r1, illegal_lockout_in, ps_stall_in}),
		.dout({leak1_i1_stall, leak1_i0_stall, dec_extint_stall, pause_state, tlu_wr_pause_r1, tlu_wr_pause_r2, illegal_lockout, ps_stall})
	);
	rvdffie #(.WIDTH(8)) misc2ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({lsu_trigger_match_m[3:0], lsu_pmu_misaligned_m, div_active_in, exu_flush_final, dec_debug_valid_d}),
		.dout({lsu_trigger_match_r[3:0], lsu_pmu_misaligned_r, div_active, flush_final_r, debug_valid_x})
	);
	generate
		if (pt[2130-:5] == 1) begin
			assign i0_brp_valid = (dec_i0_brp[50] & ~leak1_mode) & ~i0_icaf_d;
			wire [1:1] sv2v_tmp_123E1;
			assign sv2v_tmp_123E1 = 1'b0;
			always @(*) dec_i0_predict_p_d[55] = sv2v_tmp_123E1;
			wire [1:1] sv2v_tmp_D766F;
			assign sv2v_tmp_D766F = 1'b0;
			always @(*) dec_i0_predict_p_d[54] = sv2v_tmp_D766F;
			wire [1:1] sv2v_tmp_EE665;
			assign sv2v_tmp_EE665 = 1'b0;
			always @(*) dec_i0_predict_p_d[53] = sv2v_tmp_EE665;
			wire [1:1] sv2v_tmp_4A5D3;
			assign sv2v_tmp_4A5D3 = i0_pcall;
			always @(*) dec_i0_predict_p_d[34] = sv2v_tmp_4A5D3;
			wire [1:1] sv2v_tmp_C4472;
			assign sv2v_tmp_C4472 = i0_pja;
			always @(*) dec_i0_predict_p_d[33] = sv2v_tmp_C4472;
			wire [1:1] sv2v_tmp_BC36C;
			assign sv2v_tmp_BC36C = i0_pret;
			always @(*) dec_i0_predict_p_d[31] = sv2v_tmp_BC36C;
			wire [31:1] sv2v_tmp_16255;
			assign sv2v_tmp_16255 = dec_i0_brp[32:2];
			always @(*) dec_i0_predict_p_d[30:0] = sv2v_tmp_16255;
			wire [1:1] sv2v_tmp_CF546;
			assign sv2v_tmp_CF546 = dec_i0_pc4_d;
			always @(*) dec_i0_predict_p_d[52] = sv2v_tmp_CF546;
			wire [2:1] sv2v_tmp_1B1F0;
			assign sv2v_tmp_1B1F0 = dec_i0_brp[37:36];
			always @(*) dec_i0_predict_p_d[51:50] = sv2v_tmp_1B1F0;
			wire [1:1] sv2v_tmp_3FDDA;
			assign sv2v_tmp_3FDDA = i0_brp_valid & i0_legal_decode_d;
			always @(*) dec_i0_predict_p_d[37] = sv2v_tmp_3FDDA;
			assign i0_notbr_error = i0_brp_valid & ~(((i0_dp_raw[28] | i0_pcall_raw) | i0_pja_raw) | i0_pret_raw);
			assign i0_br_toffset_error = ((i0_brp_valid & dec_i0_brp[37]) & (dec_i0_brp[49:38] != i0_br_offset[11:0])) & ~i0_pret_raw;
			assign i0_ret_error = i0_brp_valid & (dec_i0_brp[0] ^ i0_pret_raw);
			assign i0_br_error = ((dec_i0_brp[35] | i0_notbr_error) | i0_br_toffset_error) | i0_ret_error;
			wire [1:1] sv2v_tmp_75A7E;
			assign sv2v_tmp_75A7E = (i0_br_error & i0_legal_decode_d) & ~leak1_mode;
			always @(*) dec_i0_predict_p_d[36] = sv2v_tmp_75A7E;
			wire [1:1] sv2v_tmp_6E7A2;
			assign sv2v_tmp_6E7A2 = (dec_i0_brp[34] & i0_legal_decode_d) & ~leak1_mode;
			always @(*) dec_i0_predict_p_d[35] = sv2v_tmp_6E7A2;
			assign i0_predict_index_d[pt[2172-:9]:pt[2163-:6]] = dec_i0_bp_index;
			assign i0_predict_btag_d[pt[2139-:9] - 1:0] = dec_i0_bp_btag[pt[2139-:9] - 1:0];
			assign i0_br_error_all = (i0_br_error | dec_i0_brp[34]) & ~leak1_mode;
			wire [12:1] sv2v_tmp_AC6BD;
			assign sv2v_tmp_AC6BD = i0_br_offset[11:0];
			always @(*) dec_i0_predict_p_d[49:38] = sv2v_tmp_AC6BD;
			assign i0_predict_fghr_d[pt[2236-:8] - 1:0] = dec_i0_bp_fghr[pt[2236-:8] - 1:0];
			wire [1:1] sv2v_tmp_11732;
			assign sv2v_tmp_11732 = dec_i0_brp[1];
			always @(*) dec_i0_predict_p_d[32] = sv2v_tmp_11732;
			if (pt[2120-:5]) begin
				wire btb_error_found;
				wire btb_error_found_f;
				wire [$clog2(pt[2061-:14]) - 1:0] fa_error_index_ns;
				assign btb_error_found = (i0_br_error_all | btb_error_found_f) & ~dec_tlu_flush_lower_r;
				assign fa_error_index_ns = (i0_br_error_all & ~btb_error_found_f ? dec_i0_bp_fa_index : dec_fa_error_index);
				rvdff #(.WIDTH($clog2(pt[2061-:14]) + 1)) btberrorfa_f(
					.rst_l(rst_l),
					.clk(active_clk),
					.din({btb_error_found, fa_error_index_ns}),
					.dout({btb_error_found_f, dec_fa_error_index})
				);
			end
			else assign dec_fa_error_index = 'b0;
		end
		else begin
			always @(*) begin
				dec_i0_predict_p_d = {56 {1'sb0}};
				dec_i0_predict_p_d[34] = i0_pcall;
				dec_i0_predict_p_d[33] = i0_pja;
				dec_i0_predict_p_d[31] = i0_pret;
				dec_i0_predict_p_d[52] = dec_i0_pc4_d;
			end
			assign i0_br_error_all = 1'b0;
			assign i0_predict_index_d = {(pt[2172-:9] >= pt[2163-:6] ? (pt[2172-:9] - pt[2163-:6]) + 1 : (pt[2163-:6] - pt[2172-:9]) + 1) {1'sb0}};
			assign i0_predict_btag_d = {pt[2139-:9] {1'sb0}};
			assign i0_predict_fghr_d = {pt[2236-:8] {1'sb0}};
			assign i0_brp_valid = 1'b0;
		end
	endgenerate
	assign i0_icaf_d = dec_i0_icaf_d | dec_i0_dbecc_d;
	assign i0_instr_error = i0_icaf_d;
	always @(*) begin
		i0_dp = i0_dp_raw;
		if (i0_br_error_all | i0_instr_error) begin
			i0_dp = {95 {1'sb0}};
			i0_dp[49] = 1'b1;
			i0_dp[48] = 1'b1;
			i0_dp[47] = 1'b1;
			i0_dp[35] = 1'b1;
			i0_dp[0] = 1'b1;
			i0_dp[13] = 1'b1;
		end
	end
	assign i0[31:0] = dec_i0_instr_d[31:0];
	assign dec_i0_select_pc_d = i0_dp[42];
	assign i0_predict_br = ((i0_dp[28] | i0_pcall) | i0_pja) | i0_pret;
	assign i0_predict_nt = ~(dec_i0_brp[37] & i0_brp_valid) & i0_predict_br;
	assign i0_predict_t = (dec_i0_brp[37] & i0_brp_valid) & i0_predict_br;
	assign i0_ap[8] = i0_dp[38];
	assign i0_ap[7] = i0_dp[37];
	assign i0_ap[18] = i0_dp[36];
	assign i0_ap[17] = i0_dp[35];
	assign i0_ap[16] = i0_dp[34];
	assign i0_ap[15] = i0_dp[33];
	assign i0_ap[14] = i0_dp[31];
	assign i0_ap[13] = i0_dp[32];
	assign i0_ap[6] = i0_dp[30];
	assign i0_ap[5] = i0_dp[29];
	assign i0_ap[12] = i0_dp[27];
	assign i0_ap[11] = i0_dp[26];
	assign i0_ap[10] = i0_dp[24];
	assign i0_ap[9] = i0_dp[25];
	assign i0_ap[43] = i0_dp[94];
	assign i0_ap[42] = i0_dp[93];
	assign i0_ap[41] = i0_dp[92];
	assign i0_ap[40] = i0_dp[91];
	assign i0_ap[39] = i0_dp[90];
	assign i0_ap[22] = i0_dp[53];
	assign i0_ap[21] = i0_dp[52];
	assign i0_ap[20] = i0_dp[51];
	assign i0_ap[19] = i0_dp[50];
	assign i0_ap[38] = i0_dp[89];
	assign i0_ap[37] = i0_dp[88];
	assign i0_ap[36] = i0_dp[87];
	assign i0_ap[35] = i0_dp[86];
	assign i0_ap[34] = i0_dp[85];
	assign i0_ap[33] = i0_dp[84];
	assign i0_ap[32] = i0_dp[83];
	assign i0_ap[31] = i0_dp[82];
	assign i0_ap[30] = i0_dp[81];
	assign i0_ap[29] = i0_dp[80];
	assign i0_ap[28] = i0_dp[79];
	assign i0_ap[27] = i0_dp[78];
	assign i0_ap[26] = i0_dp[77];
	assign i0_ap[25] = i0_dp[76];
	assign i0_ap[24] = i0_dp[75];
	assign i0_ap[23] = i0_dp[74];
	assign i0_ap[1] = i0_csr_write_only_d;
	assign i0_ap[0] = i0_dp[15];
	assign i0_ap[4] = i0_jal;
	assign i0_ap_pc2 = ~dec_i0_pc4_d;
	assign i0_ap_pc4 = dec_i0_pc4_d;
	assign i0_ap[2] = i0_predict_nt;
	assign i0_ap[3] = i0_predict_t;
	always @(*) begin
		found = 0;
		cam_wen[NBLOAD_SIZE_MSB:0] = {(NBLOAD_SIZE_MSB >= 0 ? NBLOAD_SIZE_MSB + 1 : 1 - NBLOAD_SIZE_MSB) {1'sb0}};
		begin : sv2v_autoblock_37
			reg signed [31:0] i;
			for (i = 0; i < NBLOAD_SIZE; i = i + 1)
				if (~found) begin
					if (~cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9]) begin
						cam_wen[i] = cam_write;
						found = 1'b1;
					end
					else
						cam_wen[i] = 0;
				end
				else
					cam_wen[i] = 0;
		end
	end
	assign cam_write = lsu_nonblock_load_valid_m;
	assign cam_write_tag[NBLOAD_TAG_MSB:0] = lsu_nonblock_load_tag_m[NBLOAD_TAG_MSB:0];
	assign cam_inv_reset = lsu_nonblock_load_inv_r;
	assign cam_inv_reset_tag[NBLOAD_TAG_MSB:0] = lsu_nonblock_load_inv_tag_r[NBLOAD_TAG_MSB:0];
	assign cam_data_reset = lsu_nonblock_load_data_valid | lsu_nonblock_load_data_error;
	assign cam_data_reset_tag[NBLOAD_TAG_MSB:0] = lsu_nonblock_load_data_tag[NBLOAD_TAG_MSB:0];
	assign nonblock_load_rd[4:0] = (x_d[3] ? x_d[8:4] : 5'b00000);
	generate
		genvar i;
		for (i = 0; i < NBLOAD_SIZE; i = i + 1) begin : cam_array
			assign cam_inv_reset_val[i] = (cam_inv_reset & (cam_inv_reset_tag[NBLOAD_TAG_MSB:0] == cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + ((5 + NBLOAD_TAG_MSB) >= 5 ? 5 + NBLOAD_TAG_MSB : ((5 + NBLOAD_TAG_MSB) + ((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))) - 1)-:((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))])) & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9];
			assign cam_data_reset_val[i] = (cam_data_reset & (cam_data_reset_tag[NBLOAD_TAG_MSB:0] == cam_raw[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + ((5 + NBLOAD_TAG_MSB) >= 5 ? 5 + NBLOAD_TAG_MSB : ((5 + NBLOAD_TAG_MSB) + ((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))) - 1)-:((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))])) & cam_raw[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9];
			always @(*) begin
				cam[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10] = cam_raw[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10];
				if (cam_data_reset_val[i])
					cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9] = 1'b0;
				cam_in[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10] = {10 {1'sb0}};
				if (cam_wen[i]) begin
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9] = 1'b1;
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 8] = 1'b0;
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + ((5 + NBLOAD_TAG_MSB) >= 5 ? 5 + NBLOAD_TAG_MSB : ((5 + NBLOAD_TAG_MSB) + ((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))) - 1)-:((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))] = cam_write_tag[NBLOAD_TAG_MSB:0];
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 4-:5] = nonblock_load_rd[4:0];
				end
				else if (cam_inv_reset_val[i] | ((i0_wen_r & (r_d_in[8:4] == cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 4-:5])) & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 8]))
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9] = 1'b0;
				else
					cam_in[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10] = cam[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10];
				if ((nonblock_load_valid_m_delay & (lsu_nonblock_load_inv_tag_r[NBLOAD_TAG_MSB:0] == cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + ((5 + NBLOAD_TAG_MSB) >= 5 ? 5 + NBLOAD_TAG_MSB : ((5 + NBLOAD_TAG_MSB) + ((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))) - 1)-:((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))])) & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9])
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 8] = 1'b1;
				if (dec_tlu_force_halt)
					cam_in[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9] = 1'b0;
			end
			rvdffie #(.WIDTH(10)) cam_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(cam_in[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10]),
				.dout(cam_raw[(NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10+:10])
			);
			assign nonblock_load_write[i] = (load_data_tag[NBLOAD_TAG_MSB:0] == cam_raw[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + ((5 + NBLOAD_TAG_MSB) >= 5 ? 5 + NBLOAD_TAG_MSB : ((5 + NBLOAD_TAG_MSB) + ((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))) - 1)-:((5 + NBLOAD_TAG_MSB) >= 5 ? (5 + NBLOAD_TAG_MSB) - 4 : 6 - (5 + NBLOAD_TAG_MSB))]) & cam_raw[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9];
		end
	endgenerate
	assign load_data_tag[NBLOAD_TAG_MSB:0] = lsu_nonblock_load_data_tag[NBLOAD_TAG_MSB:0];
	assign nonblock_load_cancel = (r_d_in[8:4] == dec_nonblock_load_waddr[4:0]) & i0_wen_r;
	assign dec_nonblock_load_wen = (lsu_nonblock_load_data_valid & |nonblock_load_write[NBLOAD_SIZE_MSB:0]) & ~nonblock_load_cancel;
	always @(*) begin
		dec_nonblock_load_waddr[4:0] = {5 {1'sb0}};
		i0_nonblock_load_stall = i0_nonblock_boundary_stall;
		begin : sv2v_autoblock_38
			reg signed [31:0] i;
			for (i = 0; i < NBLOAD_SIZE; i = i + 1)
				begin
					dec_nonblock_load_waddr[4:0] = dec_nonblock_load_waddr[4:0] | ({5 {nonblock_load_write[i]}} & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 4-:5]);
					i0_nonblock_load_stall = i0_nonblock_load_stall | ((dec_i0_rs1_en_d & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9]) & (cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 4-:5] == i0r[14:10]));
					i0_nonblock_load_stall = i0_nonblock_load_stall | ((dec_i0_rs2_en_d & cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 9]) & (cam[((NBLOAD_SIZE_MSB >= 0 ? i : NBLOAD_SIZE_MSB - i) * 10) + 4-:5] == i0r[9:5]));
				end
		end
	end
	assign i0_nonblock_boundary_stall = (((nonblock_load_rd[4:0] == i0r[14:10]) & lsu_nonblock_load_valid_m) & dec_i0_rs1_en_d) | (((nonblock_load_rd[4:0] == i0r[9:5]) & lsu_nonblock_load_valid_m) & dec_i0_rs2_en_d);
	rvdffs #(.WIDTH(1)) wbnbloaddelayff(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(i0_r_ctl_en),
		.din(lsu_nonblock_load_valid_m),
		.dout(nonblock_load_valid_m_delay)
	);
	assign i0_load_kill_wen_r = nonblock_load_valid_m_delay & r_d[3];
	assign csr_read = csr_ren_qual_d;
	assign csr_write = dec_csr_wen_unq_d;
	assign i0_br_unpred = i0_dp[23] & ~i0_predict_br;
	localparam [3:0] eb1_pkg_ALU = 4'b0100;
	localparam [3:0] eb1_pkg_BITMANIPU = 4'b1111;
	localparam [3:0] eb1_pkg_CONDBR = 4'b1101;
	localparam [3:0] eb1_pkg_CSRREAD = 4'b0101;
	localparam [3:0] eb1_pkg_CSRRW = 4'b0111;
	localparam [3:0] eb1_pkg_CSRWRITE = 4'b0110;
	localparam [3:0] eb1_pkg_EBREAK = 4'b1000;
	localparam [3:0] eb1_pkg_ECALL = 4'b1001;
	localparam [3:0] eb1_pkg_FENCE = 4'b1010;
	localparam [3:0] eb1_pkg_FENCEI = 4'b1011;
	localparam [3:0] eb1_pkg_JAL = 4'b1110;
	localparam [3:0] eb1_pkg_LOAD = 4'b0010;
	localparam [3:0] eb1_pkg_MRET = 4'b1100;
	localparam [3:0] eb1_pkg_MUL = 4'b0001;
	localparam [3:0] eb1_pkg_NULL = 4'b0000;
	localparam [3:0] eb1_pkg_STORE = 4'b0011;
	always @(*) begin
		i0_itype = eb1_pkg_NULL;
		if (i0_legal_decode_d) begin
			if (i0_dp[9])
				i0_itype = eb1_pkg_MUL;
			if (i0_dp[41])
				i0_itype = eb1_pkg_LOAD;
			if (i0_dp[40])
				i0_itype = eb1_pkg_STORE;
			if (i0_dp[1])
				i0_itype = eb1_pkg_ALU;
			if (((((((i0_dp[78] | i0_dp[73]) | i0_dp[70]) | i0_dp[66]) | i0_dp[63]) | i0_dp[56]) | i0_dp[54]) | i0_dp[50])
				i0_itype = eb1_pkg_BITMANIPU;
			if (csr_read & ~csr_write)
				i0_itype = eb1_pkg_CSRREAD;
			if (~csr_read & csr_write)
				i0_itype = eb1_pkg_CSRWRITE;
			if (csr_read & csr_write)
				i0_itype = eb1_pkg_CSRRW;
			if (i0_dp[12])
				i0_itype = eb1_pkg_EBREAK;
			if (i0_dp[11])
				i0_itype = eb1_pkg_ECALL;
			if (i0_dp[3])
				i0_itype = eb1_pkg_FENCE;
			if (i0_dp[2])
				i0_itype = eb1_pkg_FENCEI;
			if (i0_dp[10])
				i0_itype = eb1_pkg_MRET;
			if (i0_dp[28])
				i0_itype = eb1_pkg_CONDBR;
			if (i0_dp[23])
				i0_itype = eb1_pkg_JAL;
		end
	end
	eb1_dec_dec_ctl i0_dec(
		.inst(i0[31:0]),
		.out(i0_dp_raw)
	);
	rvdff #(.WIDTH(1)) lsu_idle_ff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din(lsu_idle_any),
		.dout(lsu_idle)
	);
	assign leak1_i1_stall_in = dec_tlu_flush_leak_one_r | (leak1_i1_stall & ~dec_tlu_flush_lower_r);
	assign leak1_mode = leak1_i1_stall;
	assign leak1_i0_stall_in = (dec_i0_decode_d & leak1_i1_stall) | (leak1_i0_stall & ~dec_tlu_flush_lower_r);
	assign i0_pcall_imm[20:1] = {i0[31], i0[19:12], i0[20], i0[30:21]};
	assign i0_pcall_12b_offset = (i0_pcall_imm[12] ? i0_pcall_imm[20:13] == 8'hff : i0_pcall_imm[20:13] == 8'h00);
	assign i0_pcall_case = (i0_pcall_12b_offset & i0_dp_raw[43]) & ((i0r[4:0] == 5'd1) | (i0r[4:0] == 5'd5));
	assign i0_pja_case = (i0_pcall_12b_offset & i0_dp_raw[43]) & ~((i0r[4:0] == 5'd1) | (i0r[4:0] == 5'd5));
	assign i0_pcall_raw = i0_dp_raw[23] & i0_pcall_case;
	assign i0_pcall = i0_dp[23] & i0_pcall_case;
	assign i0_pja_raw = i0_dp_raw[23] & i0_pja_case;
	assign i0_pja = i0_dp[23] & i0_pja_case;
	assign i0_br_offset[11:0] = (i0_pcall_raw | i0_pja_raw ? i0_pcall_imm[12:1] : {i0[31], i0[7], i0[30:25], i0[11:8]});
	assign i0_pret_case = ((i0_dp_raw[23] & i0_dp_raw[46]) & (i0r[4:0] == 5'b00000)) & ((i0r[14:10] == 5'd1) | (i0r[14:10] == 5'd5));
	assign i0_pret_raw = i0_dp_raw[23] & i0_pret_case;
	assign i0_pret = i0_dp[23] & i0_pret_case;
	assign i0_jal = ((i0_dp[23] & ~i0_pcall_case) & ~i0_pja_case) & ~i0_pret_case;
	assign dec_lsu_offset_d[11:0] = ({12 {(~dec_extint_stall & i0_dp[39]) & i0_dp[41]}} & i0[31:20]) | ({12 {(~dec_extint_stall & i0_dp[39]) & i0_dp[40]}} & {i0[31:25], i0[11:7]});
	assign div_p[2] = div_decode_d;
	assign div_p[1] = i0_dp[29];
	assign div_p[0] = i0_dp[4];
	assign mul_p[19] = mul_decode_d;
	assign mul_p[18] = i0_dp[8];
	assign mul_p[17] = i0_dp[7];
	assign mul_p[16] = i0_dp[6];
	assign mul_p[15] = i0_dp[72];
	assign mul_p[14] = i0_dp[71];
	assign mul_p[13] = i0_dp[69];
	assign mul_p[12] = i0_dp[68];
	assign mul_p[11] = i0_dp[67];
	assign mul_p[10] = i0_dp[80];
	assign mul_p[9] = i0_dp[79];
	assign mul_p[8] = i0_dp[65];
	assign mul_p[7] = i0_dp[64];
	assign mul_p[6] = i0_dp[62];
	assign mul_p[5] = i0_dp[61];
	assign mul_p[4] = i0_dp[60];
	assign mul_p[3] = i0_dp[59];
	assign mul_p[2] = i0_dp[58];
	assign mul_p[1] = i0_dp[57];
	assign mul_p[0] = i0_dp[55];
	always @(*) begin
		lsu_p = {14 {1'sb0}};
		if (dec_extint_stall) begin
			lsu_p[7] = 1'b1;
			lsu_p[9] = 1'b1;
			lsu_p[13] = 1'b1;
			lsu_p[0] = 1'b1;
		end
		else begin
			lsu_p[0] = lsu_decode_d;
			lsu_p[7] = i0_dp[41];
			lsu_p[6] = i0_dp[40];
			lsu_p[11] = i0_dp[22];
			lsu_p[10] = i0_dp[21];
			lsu_p[9] = i0_dp[20];
			lsu_p[12] = i0r[14:10] == 5'd2;
			lsu_p[2] = load_ldst_bypass_d;
			lsu_p[3] = store_data_bypass_d;
			lsu_p[1] = store_data_bypass_m;
			lsu_p[5] = i0_dp[29];
		end
	end
	assign dec_lsu_valid_raw_d = (((i0_valid_d & (i0_dp_raw[41] | i0_dp_raw[40])) & ~dma_dccm_stall_any) & ~i0_block_raw_d) | dec_extint_stall;
	assign i0r[14:10] = i0[19:15];
	assign i0r[9:5] = i0[24:20];
	assign i0r[4:0] = i0[11:7];
	assign dec_i0_rs1_en_d = i0_dp[48] & (i0r[14:10] != 5'd0);
	assign dec_i0_rs2_en_d = i0_dp[47] & (i0r[9:5] != 5'd0);
	assign i0_rd_en_d = i0_dp[45] & (i0r[4:0] != 5'd0);
	assign dec_i0_rs1_d[4:0] = i0r[14:10];
	assign dec_i0_rs2_d[4:0] = i0r[9:5];
	assign i0_jalimm20 = i0_dp[23] & i0_dp[43];
	assign i0_uiimm20 = ~i0_dp[23] & i0_dp[43];
	assign dec_csr_ren_d = i0_dp[19] & i0_valid_d;
	assign csr_ren_qual_d = i0_dp[19] & i0_legal_decode_d;
	assign csr_clr_d = i0_dp[18] & i0_legal_decode_d;
	assign csr_set_d = i0_dp[17] & i0_legal_decode_d;
	assign csr_write_d = i0_csr_write & i0_legal_decode_d;
	assign i0_csr_write_only_d = i0_csr_write & ~i0_dp[19];
	assign dec_csr_wen_unq_d = ((i0_dp[18] | i0_dp[17]) | i0_csr_write) & i0_valid_d;
	assign dec_csr_any_unq_d = any_csr_d & i0_valid_d;
	assign dec_csr_rdaddr_d[11:0] = {12 {dec_csr_any_unq_d}} & i0[31:20];
	assign dec_csr_wraddr_r[11:0] = {12 {r_d[22] & r_d[0]}} & r_d[20:9];
	assign dec_csr_wen_r = (r_d[22] & r_d[0]) & ~dec_tlu_i0_kill_writeb_r;
	assign dec_csr_stall_int_ff = ((((r_d[20:9] == 12'h300) | (r_d[20:9] == 12'h304)) & r_d[22]) & r_d[0]) & ~dec_tlu_i0_kill_writeb_wb;
	rvdff #(.WIDTH(5)) csrmiscff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din({csr_ren_qual_d, csr_clr_d, csr_set_d, csr_write_d, i0_dp[15]}),
		.dout({csr_read_x, csr_clr_x, csr_set_x, csr_write_x, csr_imm_x})
	);
	rvdffe #(.WIDTH(37)) csr_rddata_x_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_data_en & any_csr_d),
		.din({i0[19:15], dec_csr_rddata_d[31:0]}),
		.dout({csrimm_x[4:0], csr_rddata_x[31:0]})
	);
	assign csr_mask_x[31:0] = ({32 {csr_imm_x}} & {27'b000000000000000000000000000, csrimm_x[4:0]}) | ({32 {~csr_imm_x}} & exu_csr_rs1_x[31:0]);
	assign write_csr_data_x[31:0] = (({32 {csr_clr_x}} & (csr_rddata_x[31:0] & ~csr_mask_x[31:0])) | ({32 {csr_set_x}} & (csr_rddata_x[31:0] | csr_mask_x[31:0]))) | ({32 {csr_write_x}} & csr_mask_x[31:0]);
	assign clear_pause = (dec_tlu_flush_lower_r & ~dec_tlu_flush_pause_r) | (pause_state & (write_csr_data[31:1] == 31'b0000000000000000000000000000000));
	assign pause_state_in = (dec_tlu_wr_pause_r | pause_state) & ~clear_pause;
	assign dec_pause_state = pause_state;
	assign dec_pause_state_cg = (pause_state & ~tlu_wr_pause_r1) & ~tlu_wr_pause_r2;
	assign csr_data_wen = ((((csr_clr_x | csr_set_x) | csr_write_x) & csr_read_x) | dec_tlu_wr_pause_r) | pause_state;
	assign write_csr_data_in[31:0] = (pause_state ? write_csr_data[31:0] - 32'b00000000000000000000000000000001 : (dec_tlu_wr_pause_r ? dec_csr_wrdata_r[31:0] : write_csr_data_x[31:0]));
	rvdffe #(.WIDTH(32)) write_csr_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(csr_data_wen),
		.din(write_csr_data_in[31:0]),
		.dout(write_csr_data[31:0])
	);
	assign pause_stall = pause_state;
	assign dec_csr_wrdata_r[31:0] = (r_d[21] & r_d[0] ? i0_result_corr_r[31:0] : write_csr_data[31:0]);
	assign dec_i0_immed_d[31:0] = i0_immed_d[31:0];
	assign i0_immed_d[31:0] = (((({32 {i0_dp[46]}} & {{20 {i0[31]}}, i0[31:20]}) | ({32 {i0_dp[44]}} & {27'b000000000000000000000000000, i0[24:20]})) | ({32 {i0_jalimm20}} & {{12 {i0[31]}}, i0[19:12], i0[20], i0[30:21], 1'b0})) | ({32 {i0_uiimm20}} & {i0[31:12], 12'b000000000000})) | ({32 {i0_csr_write_only_d & i0_dp[15]}} & {27'b000000000000000000000000000, i0[19:15]});
	assign dec_i0_br_immed_d[12:1] = (i0_ap[2] & ~i0_dp[23] ? i0_br_offset[11:0] : {10'b0000000000, i0_ap_pc4, i0_ap_pc2});
	assign last_br_immed_d[12:1] = (i0_ap[2] ? {10'b0000000000, i0_ap_pc4, i0_ap_pc2} : i0_br_offset[11:0]);
	assign i0_valid_d = dec_ib0_valid_d;
	assign i0_load_stall_d = i0_dp[41] & (lsu_load_stall_any | dma_dccm_stall_any);
	assign i0_store_stall_d = i0_dp[40] & (lsu_store_stall_any | dma_dccm_stall_any);
	assign i0_presync = (((i0_dp[14] | dec_tlu_presync_d) | debug_fence_i) | debug_fence_raw) | dec_tlu_pipelining_disable;
	assign i0_postsync = ((i0_dp[13] | dec_tlu_postsync_d) | debug_fence_i) | (i0_csr_write_only_d & (i0[31:20] == 12'h7c2));
	assign debug_fence_i = dec_debug_fence_d & dbg_cmd_wrdata[0];
	assign debug_fence_raw = dec_debug_fence_d & dbg_cmd_wrdata[1];
	assign debug_fence = debug_fence_raw | debug_fence_i;
	assign i0_csr_write = i0_dp[16] & ~dec_debug_fence_d;
	assign presync_stall = i0_presync & prior_inflight_eff;
	assign prior_inflight_eff = (i0_dp[5] ? prior_inflight_x : prior_inflight);
	assign i0_div_prior_div_stall = i0_dp[5] & div_active;
	assign i0_block_raw_d = (((((((((((i0_dp[19] & prior_csr_write) | dec_extint_stall) | pause_stall) | leak1_i0_stall) | dec_tlu_debug_stall) | postsync_stall) | presync_stall) | ((i0_dp[3] | debug_fence) & ~lsu_idle)) | i0_nonblock_load_stall) | i0_load_block_d) | i0_nonblock_div_stall) | i0_div_prior_div_stall;
	assign i0_block_d = (i0_block_raw_d | i0_store_stall_d) | i0_load_stall_d;
	assign i0_exublock_d = i0_block_raw_d;
	assign prior_csr_write = (x_d[21] | r_d[21]) | wbd[21];
	generate
		if (pt[2207-:5] == 1) begin
			assign bitmanip_zbb_legal = 1'b1;
		end
		else assign bitmanip_zbb_legal = ~(i0_dp[78] & ~i0_dp[63]);
	endgenerate
	generate
		if (pt[2177-:5] == 1) begin
			assign bitmanip_zbs_legal = 1'b1;
		end
		else assign bitmanip_zbs_legal = ~i0_dp[73];
	endgenerate
	generate
		if (pt[2197-:5] == 1) begin
			assign bitmanip_zbe_legal = 1'b1;
		end
		else assign bitmanip_zbe_legal = ~i0_dp[70];
	endgenerate
	generate
		if (pt[2202-:5] == 1) begin
			assign bitmanip_zbc_legal = 1'b1;
		end
		else assign bitmanip_zbc_legal = ~i0_dp[66];
	endgenerate
	generate
		if (pt[2187-:5] == 1) begin
			assign bitmanip_zbp_legal = 1'b1;
		end
		else assign bitmanip_zbp_legal = ~(i0_dp[63] & ~i0_dp[78]);
	endgenerate
	generate
		if (pt[2182-:5] == 1) begin
			assign bitmanip_zbr_legal = 1'b1;
		end
		else assign bitmanip_zbr_legal = ~i0_dp[56];
	endgenerate
	generate
		if (pt[2192-:5] == 1) begin
			assign bitmanip_zbf_legal = 1'b1;
		end
		else assign bitmanip_zbf_legal = ~i0_dp[54];
	endgenerate
	generate
		if (pt[2212-:5] == 1) begin
			assign bitmanip_zba_legal = 1'b1;
		end
		else assign bitmanip_zba_legal = ~i0_dp[50];
	endgenerate
	generate
		if ((pt[2207-:5] == 1) | (pt[2187-:5] == 1)) begin
			assign bitmanip_zbb_zbp_legal = 1'b1;
		end
		else assign bitmanip_zbb_zbp_legal = ~(i0_dp[78] & i0_dp[63]);
	endgenerate
	assign any_csr_d = i0_dp[19] | i0_csr_write;
	assign bitmanip_legal = (((((((bitmanip_zbb_legal & bitmanip_zbs_legal) & bitmanip_zbe_legal) & bitmanip_zbc_legal) & bitmanip_zbp_legal) & bitmanip_zbr_legal) & bitmanip_zbf_legal) & bitmanip_zba_legal) & bitmanip_zbb_zbp_legal;
	assign i0_legal = (i0_dp[0] & (~any_csr_d | dec_csr_legal_d)) & bitmanip_legal;
	assign shift_illegal = dec_i0_decode_d & ~i0_legal;
	assign illegal_inst_en = shift_illegal & ~illegal_lockout;
	rvdffe #(.WIDTH(32)) illegal_any_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(illegal_inst_en),
		.din(i0_inst_d[31:0]),
		.dout(dec_illegal_inst[31:0])
	);
	assign illegal_lockout_in = (shift_illegal | illegal_lockout) & ~flush_final_r;
	assign dec_i0_decode_d = ((i0_valid_d & ~i0_block_d) & ~dec_tlu_flush_lower_r) & ~flush_final_r;
	assign i0_exudecode_d = ((i0_valid_d & ~i0_exublock_d) & ~dec_tlu_flush_lower_r) & ~flush_final_r;
	assign i0_legal_decode_d = dec_i0_decode_d & i0_legal;
	assign i0_exulegal_decode_d = i0_exudecode_d & i0_legal;
	assign dec_pmu_instr_decoded = dec_i0_decode_d;
	assign dec_pmu_decode_stall = i0_valid_d & ~dec_i0_decode_d;
	assign dec_pmu_postsync_stall = postsync_stall & i0_valid_d;
	assign dec_pmu_presync_stall = presync_stall & i0_valid_d;
	assign ps_stall_in = (dec_i0_decode_d & (i0_postsync | ~i0_legal)) | (ps_stall & prior_inflight_x);
	assign postsync_stall = ps_stall;
	assign prior_inflight_x = x_d[0];
	assign prior_inflight_wb = r_d[0];
	assign prior_inflight = prior_inflight_x | prior_inflight_wb;
	assign dec_i0_alu_decode_d = i0_exulegal_decode_d & i0_dp[49];
	assign dec_i0_branch_d = (i0_dp[28] | i0_dp[23]) | i0_br_error_all;
	assign lsu_decode_d = i0_legal_decode_d & i0_dp[39];
	assign mul_decode_d = i0_exulegal_decode_d & i0_dp[9];
	assign div_decode_d = i0_exulegal_decode_d & i0_dp[5];
	assign dec_qual_lsu_d = i0_dp[39];
	assign i0_rs1_depend_i0_x = (dec_i0_rs1_en_d & x_d[1]) & (x_d[8:4] == i0r[14:10]);
	assign i0_rs1_depend_i0_r = (dec_i0_rs1_en_d & r_d[1]) & (r_d[8:4] == i0r[14:10]);
	assign i0_rs2_depend_i0_x = (dec_i0_rs2_en_d & x_d[1]) & (x_d[8:4] == i0r[9:5]);
	assign i0_rs2_depend_i0_r = (dec_i0_rs2_en_d & r_d[1]) & (r_d[8:4] == i0r[9:5]);
	assign {i0_rs1_class_d, i0_rs1_depth_d[1:0]} = (i0_rs1_depend_i0_x ? {i0_x_c, 2'd1} : (i0_rs1_depend_i0_r ? {i0_r_c, 2'd2} : {5 {1'sb0}}));
	assign {i0_rs2_class_d, i0_rs2_depth_d[1:0]} = (i0_rs2_depend_i0_x ? {i0_x_c, 2'd1} : (i0_rs2_depend_i0_r ? {i0_r_c, 2'd2} : {5 {1'sb0}}));
	generate
		if (pt[202-:5] == 1) begin : genblock
			assign i0_load_block_d = (i0_rs1_class_d[1] & i0_rs1_depth_d[0]) | ((i0_rs2_class_d[1] & i0_rs2_depth_d[0]) & ~i0_dp[40]);
			assign load_ldst_bypass_d = ((i0_dp[41] | i0_dp[40]) & i0_rs1_depth_d[1]) & i0_rs1_class_d[1];
			assign store_data_bypass_d = (i0_dp[40] & i0_rs2_depth_d[1]) & i0_rs2_class_d[1];
			assign store_data_bypass_m = (i0_dp[40] & i0_rs2_depth_d[0]) & i0_rs2_class_d[1];
		end
		else begin : genblock
			assign i0_load_block_d = 1'b0;
			assign load_ldst_bypass_d = ((i0_dp[41] | i0_dp[40]) & i0_rs1_depth_d[0]) & i0_rs1_class_d[1];
			assign store_data_bypass_d = (i0_dp[40] & i0_rs2_depth_d[0]) & i0_rs2_class_d[1];
			assign store_data_bypass_m = 1'b0;
		end
	endgenerate
	assign dec_tlu_i0_valid_r = r_d[0] & ~dec_tlu_flush_lower_wb;
	assign d_t[5] = i0_legal_decode_d;
	assign d_t[16] = i0_icaf_d & i0_legal_decode_d;
	assign d_t[15] = dec_i0_icaf_second_d & i0_legal_decode_d;
	assign d_t[14:13] = dec_i0_icaf_type_d[1:0];
	assign d_t[12] = (i0_dp[2] | debug_fence_i) & i0_legal_decode_d;
	assign d_t[3-:4] = i0_itype;
	assign d_t[7] = i0_br_unpred;
	assign d_t[6] = 1'b0;
	assign d_t[4] = 1'b0;
	assign d_t[11:8] = dec_i0_trigger_match_d[3:0] & {4 {dec_i0_decode_d}};
	rvdfflie #(
		.WIDTH(17),
		.LEFT(9)
	) trap_xff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_ctl_en),
		.din(d_t),
		.dout(x_t)
	);
	always @(*) begin
		x_t_in = x_t;
		x_t_in[11:8] = x_t[11-:4] & ~{4 {dec_tlu_flush_lower_wb}};
	end
	rvdfflie #(
		.WIDTH(17),
		.LEFT(9)
	) trap_r_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_ctl_en),
		.din(x_t_in),
		.dout(r_t)
	);
	always @(*) begin
		r_t_in = r_t;
		r_t_in[11:8] = ({4 {r_d[3] | r_d[2]}} & lsu_trigger_match_r[3:0]) | r_t[11:8];
		r_t_in[4] = lsu_pmu_misaligned_r;
		if (dec_tlu_flush_lower_wb)
			r_t_in = {17 {1'sb0}};
	end
	always @(*) begin
		dec_tlu_packet_r = r_t_in;
		dec_tlu_packet_r[6] = r_d[23] & r_d[0];
	end
	assign i0_d_c[2] = i0_dp[9] & i0_legal_decode_d;
	assign i0_d_c[1] = i0_dp[41] & i0_legal_decode_d;
	assign i0_d_c[0] = i0_dp[49] & i0_legal_decode_d;
	rvdffs #(.WIDTH(3)) i0_x_c_ff(
		.rst_l(rst_l),
		.en(i0_x_ctl_en),
		.clk(active_clk),
		.din(i0_d_c),
		.dout(i0_x_c)
	);
	rvdffs #(.WIDTH(3)) i0_r_c_ff(
		.rst_l(rst_l),
		.en(i0_r_ctl_en),
		.clk(active_clk),
		.din(i0_x_c),
		.dout(i0_r_c)
	);
	assign d_d[8:4] = i0r[4:0];
	assign d_d[1] = i0_rd_en_d & i0_legal_decode_d;
	assign d_d[0] = dec_i0_decode_d;
	assign d_d[3] = i0_dp[41] & i0_legal_decode_d;
	assign d_d[2] = i0_dp[40] & i0_legal_decode_d;
	assign d_d[23] = i0_dp[5] & i0_legal_decode_d;
	assign d_d[22] = dec_csr_wen_unq_d & i0_legal_decode_d;
	assign d_d[21] = i0_csr_write_only_d & dec_i0_decode_d;
	assign d_d[20:9] = (d_d[22] ? i0[31:20] : {12 {1'sb0}});
	rvdff #(.WIDTH(3)) i0cgff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din(i0_pipe_en[3:1]),
		.dout(i0_pipe_en[2:0])
	);
	assign i0_pipe_en[3] = dec_i0_decode_d;
	assign i0_x_ctl_en = |i0_pipe_en[3:2] | clk_override;
	assign i0_r_ctl_en = |i0_pipe_en[2:1] | clk_override;
	assign i0_wb_ctl_en = |i0_pipe_en[1:0] | clk_override;
	assign i0_x_data_en = i0_pipe_en[3] | clk_override;
	assign i0_r_data_en = i0_pipe_en[2] | clk_override;
	assign i0_wb_data_en = i0_pipe_en[1] | clk_override;
	assign dec_data_en[1:0] = {i0_x_data_en, i0_r_data_en};
	assign dec_ctl_en[1:0] = {i0_x_ctl_en, i0_r_ctl_en};
	rvdfflie #(
		.WIDTH(24),
		.LEFT(15)
	) e1ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_ctl_en),
		.din(d_d),
		.dout(x_d)
	);
	always @(*) begin
		x_d_in = x_d;
		x_d_in[1] = (x_d[1] & ~dec_tlu_flush_lower_wb) & ~dec_tlu_flush_lower_r;
		x_d_in[0] = (x_d[0] & ~dec_tlu_flush_lower_wb) & ~dec_tlu_flush_lower_r;
	end
	rvdfflie #(
		.WIDTH(24),
		.LEFT(15)
	) r_d_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_r_ctl_en),
		.din(x_d_in),
		.dout(r_d)
	);
	always @(*) begin
		r_d_in = r_d;
		r_d_in[8:4] = r_d[8:4];
		r_d_in[1] = r_d[1] & ~dec_tlu_flush_lower_wb;
		r_d_in[0] = r_d[0] & ~dec_tlu_flush_lower_wb;
		r_d_in[3] = r_d[3] & ~dec_tlu_flush_lower_wb;
		r_d_in[2] = r_d[2] & ~dec_tlu_flush_lower_wb;
	end
	rvdfflie #(
		.WIDTH(24),
		.LEFT(15)
	) wbff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_wb_ctl_en),
		.din(r_d_in),
		.dout(wbd)
	);
	assign dec_i0_waddr_r[4:0] = r_d_in[8:4];
	assign i0_wen_r = r_d_in[1] & ~dec_tlu_i0_kill_writeb_r;
	assign dec_i0_wen_r = (i0_wen_r & ~r_d_in[23]) & ~i0_load_kill_wen_r;
	assign dec_i0_wdata_r[31:0] = i0_result_corr_r[31:0];
	assign div_e1_to_r = (x_d[23] & x_d[0]) | (r_d[23] & r_d[0]);
	assign div_active_in = i0_div_decode_d | ((div_active & ~exu_div_wren) & ~nonblock_div_cancel);
	assign dec_div_active = div_active;
	assign i0_nonblock_div_stall = ((dec_i0_rs1_en_d & div_active) & (div_waddr_wb[4:0] == i0r[14:10])) | ((dec_i0_rs2_en_d & div_active) & (div_waddr_wb[4:0] == i0r[9:5]));
	assign div_flush = (((x_d[23] & x_d[0]) & (x_d[8:4] == 5'b00000)) | ((x_d[23] & x_d[0]) & dec_tlu_flush_lower_r)) | (((r_d[23] & r_d[0]) & dec_tlu_flush_lower_r) & dec_tlu_i0_kill_writeb_r);
	assign nonblock_div_cancel = (div_active & div_flush) | (((div_active & ~div_e1_to_r) & (r_d[8:4] == div_waddr_wb[4:0])) & i0_wen_r);
	assign dec_div_cancel = nonblock_div_cancel;
	assign i0_div_decode_d = i0_legal_decode_d & i0_dp[5];
	generate
		if (pt[202-:5] == 1) begin : genblock1
			assign i0_result_x[31:0] = exu_i0_result_x[31:0];
			assign i0_result_r[31:0] = (r_d[1] & r_d[3] ? lsu_result_m[31:0] : i0_result_r_raw[31:0]);
		end
		else begin : genblock1
			assign i0_result_x[31:0] = (x_d[1] & x_d[3] ? lsu_result_m[31:0] : exu_i0_result_x[31:0]);
			assign i0_result_r[31:0] = i0_result_r_raw[31:0];
		end
	endgenerate
	rvdffe #(.WIDTH(32)) i0_result_r_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_r_data_en & ((x_d[1] | x_d[22]) | debug_valid_x)),
		.din(i0_result_x[31:0]),
		.dout(i0_result_r_raw[31:0])
	);
	assign i0_result_corr_r[31:0] = (r_d[1] & r_d[3] ? lsu_result_corr_r[31:0] : i0_result_r_raw[31:0]);
	rvdffe #(.WIDTH(12)) e1brpcff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_data_en),
		.din(last_br_immed_d[12:1]),
		.dout(last_br_immed_x[12:1])
	);
	assign i0_wb_en = i0_wb_data_en;
	assign i0_inst_wb_in[31:0] = i0_inst_r[31:0];
	assign i0_inst_d[31:0] = (dec_i0_pc4_d ? i0[31:0] : {16'b0000000000000000, ifu_i0_cinst[15:0]});
	assign trace_enable = ~dec_tlu_trace_disable;
	rvdffe #(
		.WIDTH(5),
		.OVERRIDE(1)
	) i0rdff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_div_decode_d),
		.din(i0r[4:0]),
		.dout(div_waddr_wb[4:0])
	);
	rvdffe #(.WIDTH(32)) i0xinstff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_x_data_en & trace_enable),
		.din(i0_inst_d[31:0]),
		.dout(i0_inst_x[31:0])
	);
	rvdffe #(.WIDTH(32)) i0cinstff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_r_data_en & trace_enable),
		.din(i0_inst_x[31:0]),
		.dout(i0_inst_r[31:0])
	);
	rvdffe #(.WIDTH(32)) i0wbinstff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_wb_en & trace_enable),
		.din(i0_inst_wb_in[31:0]),
		.dout(i0_inst_wb[31:0])
	);
	rvdffe #(.WIDTH(31)) i0wbpcff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_wb_en & trace_enable),
		.din(dec_tlu_i0_pc_r[31:1]),
		.dout(i0_pc_wb[31:1])
	);
	assign dec_i0_inst_wb[31:0] = i0_inst_wb[31:0];
	assign dec_i0_pc_wb[31:1] = i0_pc_wb[31:1];
	rvdffpcie #(.WIDTH(31)) i0_pc_r_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(i0_r_data_en),
		.din(exu_i0_pc_x[31:1]),
		.dout(dec_i0_pc_r[31:1])
	);
	assign dec_tlu_i0_pc_r[31:1] = dec_i0_pc_r[31:1];
	rvbradder ibradder_correct(
		.pc(exu_i0_pc_x[31:1]),
		.offset(last_br_immed_x[12:1]),
		.dout(pred_correct_npc_x[31:1])
	);
	assign i0_rs1_nonblock_load_bypass_en_d = (dec_i0_rs1_en_d & dec_nonblock_load_wen) & (dec_nonblock_load_waddr[4:0] == i0r[14:10]);
	assign i0_rs2_nonblock_load_bypass_en_d = (dec_i0_rs2_en_d & dec_nonblock_load_wen) & (dec_nonblock_load_waddr[4:0] == i0r[9:5]);
	assign i0_rs1bypass[2] = i0_rs1_depth_d[0] & (i0_rs1_class_d[0] | i0_rs1_class_d[2]);
	assign i0_rs1bypass[1] = i0_rs1_depth_d[0] & i0_rs1_class_d[1];
	assign i0_rs1bypass[0] = i0_rs1_depth_d[1] & ((i0_rs1_class_d[0] | i0_rs1_class_d[2]) | i0_rs1_class_d[1]);
	assign i0_rs2bypass[2] = i0_rs2_depth_d[0] & (i0_rs2_class_d[0] | i0_rs2_class_d[2]);
	assign i0_rs2bypass[1] = i0_rs2_depth_d[0] & i0_rs2_class_d[1];
	assign i0_rs2bypass[0] = i0_rs2_depth_d[1] & ((i0_rs2_class_d[0] | i0_rs2_class_d[2]) | i0_rs2_class_d[1]);
	assign dec_i0_rs1_bypass_en_d[3] = ((i0_rs1_nonblock_load_bypass_en_d & ~i0_rs1bypass[0]) & ~i0_rs1bypass[1]) & ~i0_rs1bypass[2];
	assign dec_i0_rs1_bypass_en_d[2] = i0_rs1bypass[2];
	assign dec_i0_rs1_bypass_en_d[1] = i0_rs1bypass[1];
	assign dec_i0_rs1_bypass_en_d[0] = i0_rs1bypass[0];
	assign dec_i0_rs2_bypass_en_d[3] = ((i0_rs2_nonblock_load_bypass_en_d & ~i0_rs2bypass[0]) & ~i0_rs2bypass[1]) & ~i0_rs2bypass[2];
	assign dec_i0_rs2_bypass_en_d[2] = i0_rs2bypass[2];
	assign dec_i0_rs2_bypass_en_d[1] = i0_rs2bypass[1];
	assign dec_i0_rs2_bypass_en_d[0] = i0_rs2bypass[0];
	assign dec_i0_result_r[31:0] = i0_result_r[31:0];
endmodule
module eb1_dec_dec_ctl (
	inst,
	out
);
	input wire [31:0] inst;
	output wire [94:0] out;
	wire [31:0] i;
	assign i[31:0] = inst[31:0];
	assign out[49] = (((((((((((((((((((((((i[30] & i[24]) & i[23]) & !i[22]) & !i[21]) & !i[20]) & i[14]) & !i[5]) & i[4]) | (((i[29] & !i[27]) & !i[24]) & i[4])) | (((!i[25] & !i[13]) & !i[12]) & i[4])) | (((!i[30] & !i[25]) & i[13]) & i[12])) | (((i[27] & i[25]) & i[14]) & i[4])) | (((i[29] & i[27]) & !i[14]) & i[4])) | (((i[29] & !i[14]) & i[5]) & i[4])) | (((!i[27] & !i[25]) & i[14]) & i[4])) | (((i[30] & !i[29]) & !i[13]) & i[4])) | (((!i[30] & !i[27]) & !i[25]) & i[4])) | ((i[13] & !i[5]) & i[4])) | ((!i[12] & !i[5]) & i[4])) | i[2]) | i[6]) | (((((((i[30] & i[24]) & i[23]) & i[22]) & i[21]) & i[20]) & !i[5]) & i[4])) | ((((((((!i[30] & i[29]) & !i[24]) & !i[23]) & i[22]) & i[21]) & i[20]) & !i[5]) & i[4])) | (((((((!i[30] & i[24]) & !i[23]) & !i[22]) & !i[21]) & !i[20]) & !i[5]) & i[4]);
	assign out[48] = (((((((((((((!i[14] & !i[13]) & !i[2]) | ((!i[13] & i[11]) & !i[2])) | ((i[19] & i[13]) & !i[2])) | ((!i[13] & i[10]) & !i[2])) | ((i[18] & i[13]) & !i[2])) | ((!i[13] & i[9]) & !i[2])) | ((i[17] & i[13]) & !i[2])) | ((!i[13] & i[8]) & !i[2])) | ((i[16] & i[13]) & !i[2])) | ((!i[13] & i[7]) & !i[2])) | ((i[15] & i[13]) & !i[2])) | (!i[4] & !i[3])) | (!i[6] & !i[2]);
	assign out[47] = ((i[5] & !i[4]) & !i[2]) | ((!i[6] & i[5]) & !i[2]);
	assign out[46] = ((((!i[4] & !i[3]) & i[2]) | (((i[13] & !i[5]) & i[4]) & !i[2])) | (((!i[13] & !i[12]) & i[6]) & i[4])) | (((!i[12] & !i[5]) & i[4]) & !i[2]);
	assign out[45] = ((!i[5] & !i[2]) | (i[5] & i[2])) | i[4];
	assign out[44] = ((((((i[27] & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2]) | (((((!i[30] & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((i[14] & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2]);
	assign out[43] = (i[5] & i[3]) | (i[4] & i[2]);
	assign out[42] = ((!i[5] & !i[3]) & i[2]) | (i[5] & i[3]);
	assign out[41] = (!i[5] & !i[4]) & !i[2];
	assign out[40] = (!i[6] & i[5]) & !i[4];
	assign out[39] = (!i[6] & !i[4]) & !i[2];
	assign out[38] = (((((!i[14] & !i[13]) & !i[12]) & !i[5]) & i[4]) | ((!i[5] & !i[3]) & i[2])) | (((((((!i[30] & !i[25]) & !i[14]) & !i[13]) & !i[12]) & !i[6]) & i[4]) & !i[2]);
	assign out[37] = (((((((((i[30] & !i[14]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2]) | ((((((!i[29] & !i[25]) & !i[14]) & i[13]) & !i[6]) & i[4]) & !i[2])) | (((((i[27] & i[25]) & i[14]) & !i[6]) & i[5]) & !i[2])) | ((((!i[14] & i[13]) & !i[5]) & i[4]) & !i[2])) | ((i[6] & !i[4]) & !i[2]);
	assign out[36] = ((((((!i[27] & !i[25]) & i[14]) & i[13]) & i[12]) & !i[6]) & !i[2]) | ((((i[14] & i[13]) & i[12]) & !i[5]) & !i[2]);
	assign out[35] = ((((!i[6] & i[3]) | (((((((!i[29] & !i[27]) & !i[25]) & i[14]) & i[13]) & !i[12]) & !i[6]) & !i[2])) | ((i[5] & i[4]) & i[2])) | (((!i[13] & !i[12]) & i[6]) & i[4])) | ((((i[14] & i[13]) & !i[12]) & !i[5]) & !i[2]);
	assign out[34] = (((((((!i[29] & !i[27]) & !i[25]) & i[14]) & !i[13]) & !i[12]) & i[4]) & !i[2]) | (((((i[14] & !i[13]) & !i[12]) & !i[5]) & i[4]) & !i[2]);
	assign out[33] = (((((((!i[29] & !i[27]) & !i[25]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[32] = ((((((i[30] & !i[29]) & !i[27]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[31] = ((((((((!i[30] & !i[29]) & !i[27]) & !i[25]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[30] = ((((((!i[29] & !i[25]) & !i[14]) & i[13]) & !i[6]) & i[4]) & !i[2]) | ((((!i[14] & i[13]) & !i[5]) & i[4]) & !i[2]);
	assign out[29] = ((((((((((!i[27] & i[25]) & i[14]) & i[12]) & !i[6]) & i[5]) & !i[2]) | ((((!i[14] & i[13]) & i[12]) & !i[5]) & !i[2])) | (((i[13] & i[6]) & !i[4]) & !i[2])) | ((i[14] & !i[5]) & !i[4])) | (((((!i[25] & !i[14]) & i[13]) & i[12]) & !i[6]) & !i[2])) | ((((((i[27] & i[25]) & i[14]) & i[13]) & !i[6]) & i[5]) & !i[2]);
	assign out[28] = (i[6] & !i[4]) & !i[2];
	assign out[27] = (((!i[14] & !i[12]) & i[6]) & !i[4]) & !i[2];
	assign out[26] = (((!i[14] & i[12]) & i[6]) & !i[4]) & !i[2];
	assign out[25] = (((i[14] & i[12]) & i[5]) & !i[4]) & !i[2];
	assign out[24] = (((i[14] & !i[12]) & i[5]) & !i[4]) & !i[2];
	assign out[23] = i[6] & i[2];
	assign out[22] = (((!i[13] & !i[12]) & !i[6]) & !i[4]) & !i[2];
	assign out[21] = ((i[12] & !i[6]) & !i[4]) & !i[2];
	assign out[20] = (i[13] & !i[6]) & !i[4];
	assign out[19] = ((((((i[13] & i[6]) & i[4]) | ((i[7] & i[6]) & i[4])) | ((i[8] & i[6]) & i[4])) | ((i[9] & i[6]) & i[4])) | ((i[10] & i[6]) & i[4])) | ((i[11] & i[6]) & i[4]);
	assign out[18] = (((((((i[15] & i[13]) & i[12]) & i[6]) & i[4]) | ((((i[16] & i[13]) & i[12]) & i[6]) & i[4])) | ((((i[17] & i[13]) & i[12]) & i[6]) & i[4])) | ((((i[18] & i[13]) & i[12]) & i[6]) & i[4])) | ((((i[19] & i[13]) & i[12]) & i[6]) & i[4]);
	assign out[17] = ((((((i[15] & !i[12]) & i[6]) & i[4]) | (((i[16] & !i[12]) & i[6]) & i[4])) | (((i[17] & !i[12]) & i[6]) & i[4])) | (((i[18] & !i[12]) & i[6]) & i[4])) | (((i[19] & !i[12]) & i[6]) & i[4]);
	assign out[16] = ((!i[13] & i[12]) & i[6]) & i[4];
	assign out[15] = (((((((i[14] & !i[13]) & i[6]) & i[4]) | (((i[15] & i[14]) & i[6]) & i[4])) | (((i[16] & i[14]) & i[6]) & i[4])) | (((i[17] & i[14]) & i[6]) & i[4])) | (((i[18] & i[14]) & i[6]) & i[4])) | (((i[19] & i[14]) & i[6]) & i[4]);
	assign out[14] = ((((((((((!i[5] & i[3]) | (((!i[13] & i[7]) & i[6]) & i[4])) | (((!i[13] & i[8]) & i[6]) & i[4])) | (((!i[13] & i[9]) & i[6]) & i[4])) | (((!i[13] & i[10]) & i[6]) & i[4])) | (((!i[13] & i[11]) & i[6]) & i[4])) | (((i[15] & i[13]) & i[6]) & i[4])) | (((i[16] & i[13]) & i[6]) & i[4])) | (((i[17] & i[13]) & i[6]) & i[4])) | (((i[18] & i[13]) & i[6]) & i[4])) | (((i[19] & i[13]) & i[6]) & i[4]);
	assign out[13] = ((((((((((((i[12] & !i[5]) & i[3]) | ((((!i[22] & !i[13]) & !i[12]) & i[6]) & i[4])) | (((!i[13] & i[7]) & i[6]) & i[4])) | (((!i[13] & i[8]) & i[6]) & i[4])) | (((!i[13] & i[9]) & i[6]) & i[4])) | (((!i[13] & i[10]) & i[6]) & i[4])) | (((!i[13] & i[11]) & i[6]) & i[4])) | (((i[15] & i[13]) & i[6]) & i[4])) | (((i[16] & i[13]) & i[6]) & i[4])) | (((i[17] & i[13]) & i[6]) & i[4])) | (((i[18] & i[13]) & i[6]) & i[4])) | (((i[19] & i[13]) & i[6]) & i[4]);
	assign out[12] = ((((!i[22] & i[20]) & !i[13]) & !i[12]) & i[6]) & i[4];
	assign out[11] = ((((!i[21] & !i[20]) & !i[13]) & !i[12]) & i[6]) & i[4];
	assign out[10] = (((i[29] & !i[13]) & !i[12]) & i[6]) & i[4];
	assign out[9] = (((((((((((((((((((((!i[30] & i[27]) & i[24]) & i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2]) | (((((((((i[29] & i[27]) & !i[24]) & i[23]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((((i[29] & i[27]) & !i[24]) & !i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((i[27] & !i[25]) & i[13]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((i[30] & i[27]) & i[13]) & !i[6]) & i[5]) & i[4]) & !i[2])) | (((((((((i[29] & i[27]) & i[22]) & !i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((((i[29] & i[27]) & !i[21]) & i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((((i[29] & i[27]) & !i[22]) & i[21]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((((i[30] & i[29]) & i[27]) & !i[23]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | ((((((((!i[30] & i[27]) & i[23]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | ((((((((!i[30] & !i[29]) & i[27]) & !i[25]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2])) | (((((i[25] & !i[14]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((((i[30] & !i[27]) & i[24]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((i[29] & i[27]) & i[14]) & !i[6]) & i[5]) & !i[2]);
	assign out[8] = ((((((((!i[27] & i[25]) & !i[14]) & i[13]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2]) | (((((((!i[27] & i[25]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2]);
	assign out[7] = ((((((!i[27] & i[25]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[6] = (((((i[25] & !i[14]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2];
	assign out[5] = ((((!i[27] & i[25]) & i[14]) & !i[6]) & i[5]) & !i[2];
	assign out[4] = (((((!i[27] & i[25]) & i[14]) & i[13]) & !i[6]) & i[5]) & !i[2];
	assign out[3] = !i[5] & i[3];
	assign out[2] = (i[12] & !i[5]) & i[3];
	assign out[94] = ((((((((((i[30] & !i[27]) & !i[24]) & !i[22]) & !i[21]) & !i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[93] = (((((((((i[30] & !i[27]) & !i[24]) & !i[22]) & i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[92] = ((((((((i[30] & !i[27]) & !i[24]) & i[21]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[91] = ((((((((i[30] & !i[27]) & i[22]) & !i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[90] = ((((((((i[30] & !i[27]) & i[22]) & i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[89] = (((((((!i[30] & i[29]) & !i[27]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[88] = (((((((!i[30] & i[29]) & !i[27]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[87] = (((((i[27] & i[25]) & i[14]) & !i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[86] = (((((i[27] & i[25]) & i[14]) & i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[85] = ((((((!i[30] & i[27]) & !i[25]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2];
	assign out[84] = (((((i[30] & i[27]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2];
	assign out[83] = ((((((!i[30] & i[27]) & !i[25]) & i[13]) & i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[82] = ((((((i[30] & !i[27]) & !i[14]) & i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[81] = (((((((i[30] & i[29]) & !i[27]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[78] = ((((((((((((((((((i[30] & !i[27]) & !i[24]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2]) | (((((((!i[30] & i[27]) & i[14]) & i[13]) & i[12]) & !i[6]) & i[5]) & !i[2])) | ((((((((i[30] & i[29]) & !i[27]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((i[27] & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2])) | ((((((i[30] & i[14]) & !i[13]) & !i[12]) & !i[6]) & i[5]) & !i[2])) | ((((((i[30] & !i[27]) & i[13]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((i[30] & i[29]) & !i[27]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((((((((i[30] & i[29]) & i[24]) & i[23]) & i[22]) & i[21]) & i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((((((((((!i[30] & i[29]) & i[27]) & !i[24]) & !i[23]) & i[22]) & i[21]) & i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | ((((((((((((!i[30] & i[27]) & i[24]) & !i[23]) & !i[22]) & !i[21]) & !i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | ((((((((((((i[30] & i[29]) & i[24]) & i[23]) & !i[22]) & !i[21]) & !i[20]) & i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | (((((i[27] & i[25]) & i[14]) & !i[6]) & i[5]) & !i[2]);
	assign out[77] = (((((((!i[30] & i[29]) & i[27]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[76] = ((((((i[30] & !i[29]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[75] = (((((((i[30] & i[29]) & i[27]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[74] = (((((((i[30] & !i[29]) & i[27]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[73] = (((((((i[29] & i[27]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2]) | (((((((i[30] & !i[29]) & i[27]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2]);
	assign out[72] = (((((((!i[30] & i[27]) & !i[25]) & i[13]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[71] = ((((((i[30] & i[27]) & i[13]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[70] = ((((((i[27] & !i[25]) & i[13]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[69] = ((((((i[27] & i[25]) & !i[14]) & !i[13]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[68] = (((((i[27] & !i[14]) & i[13]) & i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[67] = (((((i[27] & !i[14]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[66] = (((((i[27] & i[25]) & !i[14]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[80] = (((((((i[30] & i[29]) & i[27]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[79] = (((((((!i[30] & i[29]) & i[27]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[65] = ((((((((!i[30] & !i[29]) & i[27]) & !i[25]) & !i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[64] = ((((((((!i[30] & !i[29]) & i[27]) & !i[25]) & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2];
	assign out[63] = (((((((((((((!i[30] & i[29]) & !i[27]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2]) | (((((((!i[30] & !i[29]) & i[27]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2])) | ((((((i[30] & !i[27]) & i[13]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((i[27] & !i[25]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2])) | ((((((i[30] & i[14]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2])) | ((((((i[29] & !i[27]) & i[12]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((((!i[30] & !i[29]) & i[27]) & !i[25]) & i[12]) & !i[6]) & i[5]) & i[4]) & !i[2])) | ((((((i[29] & i[14]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[2]);
	assign out[62] = ((((((((((i[30] & !i[27]) & i[24]) & !i[23]) & !i[21]) & !i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[61] = (((((((((i[30] & !i[27]) & i[24]) & !i[23]) & i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[60] = (((((((((i[30] & !i[27]) & i[24]) & !i[23]) & i[21]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[59] = (((((((((i[30] & !i[27]) & i[23]) & !i[21]) & !i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[58] = ((((((((i[30] & !i[27]) & i[23]) & i[20]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[57] = ((((((((i[30] & !i[27]) & i[23]) & i[21]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[56] = (((((((i[30] & !i[27]) & i[24]) & !i[14]) & !i[13]) & i[12]) & !i[5]) & i[4]) & !i[2];
	assign out[55] = (((((i[30] & i[27]) & i[13]) & i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[54] = (((((i[30] & i[27]) & i[13]) & i[12]) & !i[6]) & i[5]) & !i[2];
	assign out[53] = (((((i[29] & !i[14]) & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[52] = (((((i[29] & i[14]) & !i[13]) & !i[12]) & i[5]) & i[4]) & !i[2];
	assign out[51] = ((((i[29] & i[14]) & i[13]) & !i[6]) & i[5]) & !i[2];
	assign out[50] = ((((i[29] & !i[12]) & !i[6]) & i[5]) & i[4]) & !i[2];
	assign out[1] = (((((((((i[28] & i[22]) & !i[13]) & !i[12]) & i[4]) | (((((!i[30] & !i[29]) & !i[27]) & !i[25]) & !i[6]) & i[4])) | ((((((!i[29] & !i[27]) & !i[25]) & !i[13]) & i[12]) & !i[6]) & i[4])) | (((((!i[29] & !i[27]) & !i[25]) & !i[14]) & !i[6]) & i[4])) | ((i[13] & !i[5]) & i[4])) | (i[4] & i[2])) | ((!i[12] & !i[5]) & i[4]);
	assign out[0] = (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((!i[31] & !i[30]) & !i[29]) & i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[24]) & !i[23]) & i[22]) & !i[21]) & i[20]) & !i[19]) & !i[18]) & !i[17]) & !i[16]) & !i[15]) & !i[14]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & i[6]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0]) | (((((((((((((((((((((((((((((!i[31] & !i[30]) & i[29]) & i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[24]) & !i[23]) & !i[22]) & i[21]) & !i[20]) & !i[19]) & !i[18]) & !i[17]) & !i[16]) & !i[15]) & !i[14]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & i[6]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((((((((((((((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[24]) & !i[23]) & !i[22]) & !i[21]) & !i[19]) & !i[18]) & !i[17]) & !i[16]) & !i[15]) & !i[14]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((((((((!i[31] & i[29]) & !i[28]) & !i[26]) & !i[25]) & i[24]) & !i[22]) & !i[20]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((((!i[31] & i[29]) & !i[28]) & !i[26]) & !i[25]) & i[24]) & !i[22]) & !i[21]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((((!i[31] & i[29]) & !i[28]) & !i[26]) & !i[25]) & !i[23]) & !i[22]) & !i[20]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((((!i[31] & i[29]) & !i[28]) & !i[26]) & !i[25]) & !i[24]) & !i[23]) & !i[21]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[26]) & i[25]) & i[13]) & !i[6]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[30]) & !i[28]) & !i[26]) & !i[25]) & !i[24]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & !i[30]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & i[14]) & !i[12]) & !i[6]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & !i[30]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & i[13]) & !i[12]) & !i[6]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & !i[29]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[13]) & !i[12]) & !i[6]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[28]) & !i[27]) & !i[26]) & !i[25]) & i[14]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[26]) & !i[13]) & i[12]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[26]) & i[14]) & !i[6]) & i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & i[30]) & !i[28]) & i[27]) & !i[26]) & !i[25]) & !i[13]) & i[12]) & !i[6]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & i[29]) & !i[28]) & i[27]) & !i[26]) & !i[25]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[30]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[27]) & !i[26]) & !i[6]) & i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((!i[14] & !i[13]) & !i[12]) & i[6]) & i[5]) & !i[4]) & !i[3]) & i[1]) & i[0])) | (((((((((((!i[31] & !i[29]) & !i[28]) & !i[26]) & !i[25]) & i[14]) & !i[6]) & i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | ((((((((((((!i[31] & i[29]) & !i[28]) & !i[26]) & !i[25]) & !i[13]) & i[12]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((i[14] & i[6]) & i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((!i[14] & !i[13]) & i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | ((((((!i[12] & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((((!i[13] & i[12]) & i[6]) & i[5]) & !i[3]) & !i[2]) & i[1]) & i[0])) | ((((((((((((((((((((((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[27]) & !i[26]) & !i[25]) & !i[24]) & !i[23]) & !i[22]) & !i[21]) & !i[20]) & !i[19]) & !i[18]) & !i[17]) & !i[16]) & !i[15]) & !i[14]) & !i[13]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & !i[6]) & !i[5]) & !i[4]) & i[3]) & i[2]) & i[1]) & i[0])) | (((((((((((((((((((((((!i[31] & !i[30]) & !i[29]) & !i[28]) & !i[19]) & !i[18]) & !i[17]) & !i[16]) & !i[15]) & !i[14]) & !i[13]) & !i[12]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & !i[6]) & !i[5]) & !i[4]) & i[3]) & i[2]) & i[1]) & i[0])) | (((((((i[13] & i[6]) & i[5]) & i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | ((((((i[6] & i[5]) & !i[4]) & i[3]) & i[2]) & i[1]) & i[0])) | (((((((!i[14] & !i[12]) & !i[6]) & !i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | (((((((!i[13] & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1]) & i[0])) | ((((((i[13] & !i[6]) & !i[5]) & i[4]) & !i[3]) & i[1]) & i[0])) | (((((!i[6] & i[4]) & !i[3]) & i[2]) & i[1]) & i[0]);
endmodule
module eb1_dec_gpr_ctl (
	raddr0,
	raddr1,
	wen0,
	waddr0,
	wd0,
	wen1,
	waddr1,
	wd1,
	wen2,
	waddr2,
	wd2,
	clk,
	rst_l,
	rd0,
	rd1,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [4:0] raddr0;
	input wire [4:0] raddr1;
	input wire wen0;
	input wire [4:0] waddr0;
	input wire [31:0] wd0;
	input wire wen1;
	input wire [4:0] waddr1;
	input wire [31:0] wd1;
	input wire wen2;
	input wire [4:0] waddr2;
	input wire [31:0] wd2;
	input wire clk;
	input wire rst_l;
	output reg [31:0] rd0;
	output reg [31:0] rd1;
	input wire scan_mode;
	wire [1023:32] gpr_out;
	reg [1023:32] gpr_in;
	reg [31:1] w0v;
	reg [31:1] w1v;
	reg [31:1] w2v;
	wire [31:1] gpr_wr_en;
	assign gpr_wr_en[31:1] = (w0v[31:1] | w1v[31:1]) | w2v[31:1];
	generate
		genvar j;
		for (j = 1; j < 32; j = j + 1) begin : gpr
			rvdffe #(.WIDTH(32)) gprff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(gpr_wr_en[j]),
				.din(gpr_in[(j * 32) + 31-:32]),
				.dout(gpr_out[(j * 32) + 31-:32])
			);
		end
	endgenerate
	function automatic signed [4:0] sv2v_cast_5_signed;
		input reg signed [4:0] inp;
		sv2v_cast_5_signed = inp;
	endfunction
	always @(*) begin
		rd0[31:0] = 32'b00000000000000000000000000000000;
		rd1[31:0] = 32'b00000000000000000000000000000000;
		w0v[31:1] = 31'b0000000000000000000000000000000;
		w1v[31:1] = 31'b0000000000000000000000000000000;
		w2v[31:1] = 31'b0000000000000000000000000000000;
		gpr_in[32+:992] = {992 {1'sb0}};
		begin : sv2v_autoblock_39
			reg signed [31:0] j;
			for (j = 1; j < 32; j = j + 1)
				begin
					rd0[31:0] = rd0[31:0] | ({32 {raddr0[4:0] == sv2v_cast_5_signed(j)}} & gpr_out[(j * 32) + 31-:32]);
					rd1[31:0] = rd1[31:0] | ({32 {raddr1[4:0] == sv2v_cast_5_signed(j)}} & gpr_out[(j * 32) + 31-:32]);
				end
		end
		begin : sv2v_autoblock_40
			reg signed [31:0] j;
			for (j = 1; j < 32; j = j + 1)
				begin
					w0v[j] = wen0 & (waddr0[4:0] == sv2v_cast_5_signed(j));
					w1v[j] = wen1 & (waddr1[4:0] == sv2v_cast_5_signed(j));
					w2v[j] = wen2 & (waddr2[4:0] == sv2v_cast_5_signed(j));
					gpr_in[j * 32+:32] = (({32 {w0v[j]}} & wd0[31:0]) | ({32 {w1v[j]}} & wd1[31:0])) | ({32 {w2v[j]}} & wd2[31:0]);
				end
		end
	end
endmodule
module eb1_dec_ib_ctl (
	dbg_cmd_valid,
	dbg_cmd_write,
	dbg_cmd_type,
	dbg_cmd_addr,
	i0_brp,
	ifu_i0_bp_index,
	ifu_i0_bp_fghr,
	ifu_i0_bp_btag,
	ifu_i0_fa_index,
	ifu_i0_pc4,
	ifu_i0_valid,
	ifu_i0_icaf,
	ifu_i0_icaf_type,
	ifu_i0_icaf_second,
	ifu_i0_dbecc,
	ifu_i0_instr,
	ifu_i0_pc,
	dec_ib0_valid_d,
	dec_debug_valid_d,
	dec_i0_instr_d,
	dec_i0_pc_d,
	dec_i0_pc4_d,
	dec_i0_brp,
	dec_i0_bp_index,
	dec_i0_bp_fghr,
	dec_i0_bp_btag,
	dec_i0_bp_fa_index,
	dec_i0_icaf_d,
	dec_i0_icaf_second_d,
	dec_i0_icaf_type_d,
	dec_i0_dbecc_d,
	dec_debug_wdata_rs1_d,
	dec_debug_fence_d
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire dbg_cmd_valid;
	input wire dbg_cmd_write;
	input wire [1:0] dbg_cmd_type;
	input wire [31:0] dbg_cmd_addr;
	input wire [50:0] i0_brp;
	input wire [pt[2172-:9]:pt[2163-:6]] ifu_i0_bp_index;
	input wire [pt[2236-:8] - 1:0] ifu_i0_bp_fghr;
	input wire [pt[2139-:9] - 1:0] ifu_i0_bp_btag;
	input wire [$clog2(pt[2061-:14]) - 1:0] ifu_i0_fa_index;
	input wire ifu_i0_pc4;
	input wire ifu_i0_valid;
	input wire ifu_i0_icaf;
	input wire [1:0] ifu_i0_icaf_type;
	input wire ifu_i0_icaf_second;
	input wire ifu_i0_dbecc;
	input wire [31:0] ifu_i0_instr;
	input wire [31:1] ifu_i0_pc;
	output wire dec_ib0_valid_d;
	output wire dec_debug_valid_d;
	output wire [31:0] dec_i0_instr_d;
	output wire [31:1] dec_i0_pc_d;
	output wire dec_i0_pc4_d;
	output wire [50:0] dec_i0_brp;
	output wire [pt[2172-:9]:pt[2163-:6]] dec_i0_bp_index;
	output wire [pt[2236-:8] - 1:0] dec_i0_bp_fghr;
	output wire [pt[2139-:9] - 1:0] dec_i0_bp_btag;
	output wire [$clog2(pt[2061-:14]) - 1:0] dec_i0_bp_fa_index;
	output wire dec_i0_icaf_d;
	output wire dec_i0_icaf_second_d;
	output wire [1:0] dec_i0_icaf_type_d;
	output wire dec_i0_dbecc_d;
	output wire dec_debug_wdata_rs1_d;
	output wire dec_debug_fence_d;
	wire debug_valid;
	wire [4:0] dreg;
	wire [11:0] dcsr;
	wire [31:0] ib0;
	wire [31:0] ib0_debug_in;
	wire debug_read;
	wire debug_write;
	wire debug_read_gpr;
	wire debug_write_gpr;
	wire debug_read_csr;
	wire debug_write_csr;
	wire [34:0] ifu_i0_pcdata;
	wire [34:0] pc0;
	assign ifu_i0_pcdata[34:0] = {ifu_i0_icaf_second, ifu_i0_dbecc, ifu_i0_icaf, ifu_i0_pc[31:1], ifu_i0_pc4};
	assign pc0[34:0] = ifu_i0_pcdata[34:0];
	assign dec_i0_icaf_second_d = pc0[34];
	assign dec_i0_dbecc_d = pc0[33];
	assign dec_i0_icaf_d = pc0[32];
	assign dec_i0_pc_d[31:1] = pc0[31:1];
	assign dec_i0_pc4_d = pc0[0];
	assign dec_i0_icaf_type_d[1:0] = ifu_i0_icaf_type[1:0];
	assign debug_valid = dbg_cmd_valid & (dbg_cmd_type[1:0] != 2'h2);
	assign debug_read = debug_valid & ~dbg_cmd_write;
	assign debug_write = debug_valid & dbg_cmd_write;
	assign debug_read_gpr = debug_read & (dbg_cmd_type[1:0] == 2'h0);
	assign debug_write_gpr = debug_write & (dbg_cmd_type[1:0] == 2'h0);
	assign debug_read_csr = debug_read & (dbg_cmd_type[1:0] == 2'h1);
	assign debug_write_csr = debug_write & (dbg_cmd_type[1:0] == 2'h1);
	assign dreg[4:0] = dbg_cmd_addr[4:0];
	assign dcsr[11:0] = dbg_cmd_addr[11:0];
	assign ib0_debug_in[31:0] = ((({32 {debug_read_gpr}} & {12'b000000000000, dreg[4:0], 15'b110000000110011}) | ({32 {debug_write_gpr}} & {20'b00000000000000000110, dreg[4:0], 7'b0110011})) | ({32 {debug_read_csr}} & {dcsr[11:0], 20'b00000010000001110011})) | ({32 {debug_write_csr}} & {dcsr[11:0], 20'b00000001000001110011});
	assign dec_debug_wdata_rs1_d = debug_write_gpr | debug_write_csr;
	assign dec_debug_fence_d = debug_write_csr & (dcsr[11:0] == 12'h7c4);
	assign ib0[31:0] = (debug_valid ? ib0_debug_in[31:0] : ifu_i0_instr[31:0]);
	assign dec_ib0_valid_d = ifu_i0_valid | debug_valid;
	assign dec_debug_valid_d = debug_valid;
	assign dec_i0_instr_d[31:0] = ib0[31:0];
	assign dec_i0_brp = i0_brp;
	assign dec_i0_bp_index = ifu_i0_bp_index;
	assign dec_i0_bp_fghr = ifu_i0_bp_fghr;
	assign dec_i0_bp_btag = ifu_i0_bp_btag;
	assign dec_i0_bp_fa_index = ifu_i0_fa_index;
endmodule
module eb1_dec_tlu_ctl (
	clk,
	free_clk,
	free_l2clk,
	rst_l,
	scan_mode,
	rst_vec,
	nmi_int,
	nmi_vec,
	i_cpu_halt_req,
	i_cpu_run_req,
	lsu_fastint_stall_any,
	ifu_pmu_instr_aligned,
	ifu_pmu_fetch_stall,
	ifu_pmu_ic_miss,
	ifu_pmu_ic_hit,
	ifu_pmu_bus_error,
	ifu_pmu_bus_busy,
	ifu_pmu_bus_trxn,
	dec_pmu_instr_decoded,
	dec_pmu_decode_stall,
	dec_pmu_presync_stall,
	dec_pmu_postsync_stall,
	lsu_store_stall_any,
	dma_dccm_stall_any,
	dma_iccm_stall_any,
	exu_pmu_i0_br_misp,
	exu_pmu_i0_br_ataken,
	exu_pmu_i0_pc4,
	lsu_pmu_bus_trxn,
	lsu_pmu_bus_misaligned,
	lsu_pmu_bus_error,
	lsu_pmu_bus_busy,
	lsu_pmu_load_external_m,
	lsu_pmu_store_external_m,
	dma_pmu_dccm_read,
	dma_pmu_dccm_write,
	dma_pmu_any_read,
	dma_pmu_any_write,
	lsu_fir_addr,
	lsu_fir_error,
	iccm_dma_sb_error,
	lsu_error_pkt_r,
	lsu_single_ecc_error_incr,
	dec_pause_state,
	lsu_imprecise_error_store_any,
	lsu_imprecise_error_load_any,
	lsu_imprecise_error_addr_any,
	dec_csr_wen_unq_d,
	dec_csr_any_unq_d,
	dec_csr_rdaddr_d,
	dec_csr_wen_r,
	dec_csr_wraddr_r,
	dec_csr_wrdata_r,
	dec_csr_stall_int_ff,
	dec_tlu_i0_valid_r,
	exu_npc_r,
	dec_tlu_i0_pc_r,
	dec_tlu_packet_r,
	dec_illegal_inst,
	dec_i0_decode_d,
	exu_i0_br_hist_r,
	exu_i0_br_error_r,
	exu_i0_br_start_error_r,
	exu_i0_br_valid_r,
	exu_i0_br_mp_r,
	exu_i0_br_middle_r,
	exu_i0_br_way_r,
	dec_tlu_core_empty,
	dec_dbg_cmd_done,
	dec_dbg_cmd_fail,
	dec_tlu_dbg_halted,
	dec_tlu_debug_mode,
	dec_tlu_resume_ack,
	dec_tlu_debug_stall,
	dec_tlu_flush_noredir_r,
	dec_tlu_mpc_halted_only,
	dec_tlu_flush_leak_one_r,
	dec_tlu_flush_err_r,
	dec_tlu_flush_extint,
	dec_tlu_meihap,
	dbg_halt_req,
	dbg_resume_req,
	ifu_miss_state_idle,
	lsu_idle_any,
	dec_div_active,
	trigger_pkt_any,
	ifu_ic_error_start,
	ifu_iccm_rd_ecc_single_err,
	ifu_ic_debug_rd_data,
	ifu_ic_debug_rd_data_valid,
	dec_tlu_ic_diag_pkt,
	pic_claimid,
	pic_pl,
	mhwakeup,
	mexintpend,
	timer_int,
	soft_int,
	o_cpu_halt_status,
	o_cpu_halt_ack,
	o_cpu_run_ack,
	o_debug_mode_status,
	core_id,
	mpc_debug_halt_req,
	mpc_debug_run_req,
	mpc_reset_run_req,
	mpc_debug_halt_ack,
	mpc_debug_run_ack,
	debug_brkpt_status,
	dec_tlu_meicurpl,
	dec_tlu_meipt,
	dec_csr_rddata_d,
	dec_csr_legal_d,
	dec_tlu_br0_r_pkt,
	dec_tlu_i0_kill_writeb_wb,
	dec_tlu_flush_lower_wb,
	dec_tlu_i0_commit_cmt,
	dec_tlu_i0_kill_writeb_r,
	dec_tlu_flush_lower_r,
	dec_tlu_flush_path_r,
	dec_tlu_fence_i_r,
	dec_tlu_wr_pause_r,
	dec_tlu_flush_pause_r,
	dec_tlu_presync_d,
	dec_tlu_postsync_d,
	dec_tlu_mrac_ff,
	dec_tlu_force_halt,
	dec_tlu_perfcnt0,
	dec_tlu_perfcnt1,
	dec_tlu_perfcnt2,
	dec_tlu_perfcnt3,
	dec_tlu_i0_exc_valid_wb1,
	dec_tlu_i0_valid_wb1,
	dec_tlu_int_valid_wb1,
	dec_tlu_exc_cause_wb1,
	dec_tlu_mtval_wb1,
	dec_tlu_external_ldfwd_disable,
	dec_tlu_sideeffect_posted_disable,
	dec_tlu_core_ecc_disable,
	dec_tlu_bpred_disable,
	dec_tlu_wb_coalescing_disable,
	dec_tlu_pipelining_disable,
	dec_tlu_trace_disable,
	dec_tlu_dma_qos_prty,
	dec_tlu_misc_clk_override,
	dec_tlu_dec_clk_override,
	dec_tlu_ifu_clk_override,
	dec_tlu_lsu_clk_override,
	dec_tlu_bus_clk_override,
	dec_tlu_pic_clk_override,
	dec_tlu_picio_clk_override,
	dec_tlu_dccm_clk_override,
	dec_tlu_icm_clk_override
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire free_clk;
	input wire free_l2clk;
	input wire rst_l;
	input wire scan_mode;
	input wire [31:1] rst_vec;
	input wire nmi_int;
	input wire [31:1] nmi_vec;
	input wire i_cpu_halt_req;
	input wire i_cpu_run_req;
	input wire lsu_fastint_stall_any;
	input wire ifu_pmu_instr_aligned;
	input wire ifu_pmu_fetch_stall;
	input wire ifu_pmu_ic_miss;
	input wire ifu_pmu_ic_hit;
	input wire ifu_pmu_bus_error;
	input wire ifu_pmu_bus_busy;
	input wire ifu_pmu_bus_trxn;
	input wire dec_pmu_instr_decoded;
	input wire dec_pmu_decode_stall;
	input wire dec_pmu_presync_stall;
	input wire dec_pmu_postsync_stall;
	input wire lsu_store_stall_any;
	input wire dma_dccm_stall_any;
	input wire dma_iccm_stall_any;
	input wire exu_pmu_i0_br_misp;
	input wire exu_pmu_i0_br_ataken;
	input wire exu_pmu_i0_pc4;
	input wire lsu_pmu_bus_trxn;
	input wire lsu_pmu_bus_misaligned;
	input wire lsu_pmu_bus_error;
	input wire lsu_pmu_bus_busy;
	input wire lsu_pmu_load_external_m;
	input wire lsu_pmu_store_external_m;
	input wire dma_pmu_dccm_read;
	input wire dma_pmu_dccm_write;
	input wire dma_pmu_any_read;
	input wire dma_pmu_any_write;
	input wire [31:1] lsu_fir_addr;
	input wire [1:0] lsu_fir_error;
	input wire iccm_dma_sb_error;
	input wire [39:0] lsu_error_pkt_r;
	input wire lsu_single_ecc_error_incr;
	input wire dec_pause_state;
	input wire lsu_imprecise_error_store_any;
	input wire lsu_imprecise_error_load_any;
	input wire [31:0] lsu_imprecise_error_addr_any;
	input wire dec_csr_wen_unq_d;
	input wire dec_csr_any_unq_d;
	input wire [11:0] dec_csr_rdaddr_d;
	input wire dec_csr_wen_r;
	input wire [11:0] dec_csr_wraddr_r;
	input wire [31:0] dec_csr_wrdata_r;
	input wire dec_csr_stall_int_ff;
	input wire dec_tlu_i0_valid_r;
	input wire [31:1] exu_npc_r;
	input wire [31:1] dec_tlu_i0_pc_r;
	input wire [16:0] dec_tlu_packet_r;
	input wire [31:0] dec_illegal_inst;
	input wire dec_i0_decode_d;
	input wire [1:0] exu_i0_br_hist_r;
	input wire exu_i0_br_error_r;
	input wire exu_i0_br_start_error_r;
	input wire exu_i0_br_valid_r;
	input wire exu_i0_br_mp_r;
	input wire exu_i0_br_middle_r;
	input wire exu_i0_br_way_r;
	output wire dec_tlu_core_empty;
	output wire dec_dbg_cmd_done;
	output wire dec_dbg_cmd_fail;
	output wire dec_tlu_dbg_halted;
	output wire dec_tlu_debug_mode;
	output wire dec_tlu_resume_ack;
	output wire dec_tlu_debug_stall;
	output wire dec_tlu_flush_noredir_r;
	output wire dec_tlu_mpc_halted_only;
	output wire dec_tlu_flush_leak_one_r;
	output wire dec_tlu_flush_err_r;
	output wire dec_tlu_flush_extint;
	output wire [31:2] dec_tlu_meihap;
	input wire dbg_halt_req;
	input wire dbg_resume_req;
	input wire ifu_miss_state_idle;
	input wire lsu_idle_any;
	input wire dec_div_active;
	output wire [151:0] trigger_pkt_any;
	input wire ifu_ic_error_start;
	input wire ifu_iccm_rd_ecc_single_err;
	input wire [70:0] ifu_ic_debug_rd_data;
	input wire ifu_ic_debug_rd_data_valid;
	output wire [89:0] dec_tlu_ic_diag_pkt;
	input wire [7:0] pic_claimid;
	input wire [3:0] pic_pl;
	input wire mhwakeup;
	input wire mexintpend;
	input wire timer_int;
	input wire soft_int;
	output wire o_cpu_halt_status;
	output wire o_cpu_halt_ack;
	output wire o_cpu_run_ack;
	output wire o_debug_mode_status;
	input wire [31:4] core_id;
	input wire mpc_debug_halt_req;
	input wire mpc_debug_run_req;
	input wire mpc_reset_run_req;
	output wire mpc_debug_halt_ack;
	output wire mpc_debug_run_ack;
	output wire debug_brkpt_status;
	output wire [3:0] dec_tlu_meicurpl;
	output wire [3:0] dec_tlu_meipt;
	output wire [31:0] dec_csr_rddata_d;
	output wire dec_csr_legal_d;
	output wire [6:0] dec_tlu_br0_r_pkt;
	output wire dec_tlu_i0_kill_writeb_wb;
	output wire dec_tlu_flush_lower_wb;
	output wire dec_tlu_i0_commit_cmt;
	output wire dec_tlu_i0_kill_writeb_r;
	output wire dec_tlu_flush_lower_r;
	output wire [31:1] dec_tlu_flush_path_r;
	output wire dec_tlu_fence_i_r;
	output wire dec_tlu_wr_pause_r;
	output wire dec_tlu_flush_pause_r;
	output wire dec_tlu_presync_d;
	output wire dec_tlu_postsync_d;
	output wire [31:0] dec_tlu_mrac_ff;
	output wire dec_tlu_force_halt;
	output wire dec_tlu_perfcnt0;
	output wire dec_tlu_perfcnt1;
	output wire dec_tlu_perfcnt2;
	output wire dec_tlu_perfcnt3;
	output wire dec_tlu_i0_exc_valid_wb1;
	output wire dec_tlu_i0_valid_wb1;
	output wire dec_tlu_int_valid_wb1;
	output wire [4:0] dec_tlu_exc_cause_wb1;
	output wire [31:0] dec_tlu_mtval_wb1;
	output wire dec_tlu_external_ldfwd_disable;
	output wire dec_tlu_sideeffect_posted_disable;
	output wire dec_tlu_core_ecc_disable;
	output wire dec_tlu_bpred_disable;
	output wire dec_tlu_wb_coalescing_disable;
	output wire dec_tlu_pipelining_disable;
	output wire dec_tlu_trace_disable;
	output wire [2:0] dec_tlu_dma_qos_prty;
	output wire dec_tlu_misc_clk_override;
	output wire dec_tlu_dec_clk_override;
	output wire dec_tlu_ifu_clk_override;
	output wire dec_tlu_lsu_clk_override;
	output wire dec_tlu_bus_clk_override;
	output wire dec_tlu_pic_clk_override;
	output wire dec_tlu_picio_clk_override;
	output wire dec_tlu_dccm_clk_override;
	output wire dec_tlu_icm_clk_override;
	wire clk_override;
	wire e4e5_int_clk;
	wire nmi_fir_type;
	wire nmi_lsu_load_type;
	wire nmi_lsu_store_type;
	wire nmi_int_detected_f;
	wire nmi_lsu_load_type_f;
	wire nmi_lsu_store_type_f;
	wire allow_dbg_halt_csr_write;
	wire dbg_cmd_done_ns;
	wire i_cpu_run_req_d1_raw;
	wire debug_mode_status;
	wire lsu_single_ecc_error_r_d1;
	wire sel_npc_r;
	wire sel_npc_resume;
	wire ce_int;
	wire nmi_in_debug_mode;
	wire dpc_capture_npc;
	wire dpc_capture_pc;
	wire tdata_load;
	wire tdata_opcode;
	wire tdata_action;
	wire perfcnt_halted;
	wire tdata_chain;
	wire tdata_kill_write;
	wire reset_delayed;
	wire reset_detect;
	wire reset_detected;
	wire wr_mstatus_r;
	wire wr_mtvec_r;
	wire wr_mcyclel_r;
	wire wr_mcycleh_r;
	wire wr_minstretl_r;
	wire wr_minstreth_r;
	wire wr_mscratch_r;
	wire wr_mepc_r;
	wire wr_mcause_r;
	wire wr_mscause_r;
	wire wr_mtval_r;
	wire wr_mrac_r;
	wire wr_meihap_r;
	wire wr_meicurpl_r;
	wire wr_meipt_r;
	wire wr_dcsr_r;
	wire wr_dpc_r;
	wire wr_meicidpl_r;
	wire wr_meivt_r;
	wire wr_meicpct_r;
	wire wr_micect_r;
	wire wr_miccmect_r;
	wire wr_mfdht_r;
	wire wr_mfdhs_r;
	wire wr_mdccmect_r;
	wire wr_mhpme3_r;
	wire wr_mhpme4_r;
	wire wr_mhpme5_r;
	wire wr_mhpme6_r;
	wire wr_mpmc_r;
	wire [1:1] mpmc_b_ns;
	wire [1:1] mpmc;
	wire [1:1] mpmc_b;
	wire set_mie_pmu_fw_halt;
	wire fw_halted_ns;
	wire fw_halted;
	wire wr_mcountinhibit_r;
	wire [6:0] mcountinhibit;
	wire wr_mtsel_r;
	wire wr_mtdata1_t0_r;
	wire wr_mtdata1_t1_r;
	wire wr_mtdata1_t2_r;
	wire wr_mtdata1_t3_r;
	wire wr_mtdata2_t0_r;
	wire wr_mtdata2_t1_r;
	wire wr_mtdata2_t2_r;
	wire wr_mtdata2_t3_r;
	wire [31:0] mtdata2_t0;
	wire [31:0] mtdata2_t1;
	wire [31:0] mtdata2_t2;
	wire [31:0] mtdata2_t3;
	wire [31:0] mtdata2_tsel_out;
	wire [31:0] mtdata1_tsel_out;
	wire [9:0] mtdata1_t0_ns;
	wire [9:0] mtdata1_t0;
	wire [9:0] mtdata1_t1_ns;
	wire [9:0] mtdata1_t1;
	wire [9:0] mtdata1_t2_ns;
	wire [9:0] mtdata1_t2;
	wire [9:0] mtdata1_t3_ns;
	wire [9:0] mtdata1_t3;
	wire [9:0] tdata_wrdata_r;
	wire [1:0] mtsel_ns;
	wire [1:0] mtsel;
	wire tlu_i0_kill_writeb_r;
	wire [1:0] mstatus_ns;
	wire [1:0] mstatus;
	wire [1:0] mfdhs_ns;
	wire [1:0] mfdhs;
	wire [31:0] force_halt_ctr;
	wire [31:0] force_halt_ctr_f;
	wire force_halt;
	wire [5:0] mfdht;
	wire [5:0] mfdht_ns;
	wire mstatus_mie_ns;
	wire [30:0] mtvec_ns;
	wire [30:0] mtvec;
	wire [15:2] dcsr_ns;
	wire [15:2] dcsr;
	wire [5:0] mip_ns;
	wire [5:0] mip;
	wire [5:0] mie_ns;
	wire [5:0] mie;
	wire [31:0] mcyclel_ns;
	wire [31:0] mcyclel;
	wire [31:0] mcycleh_ns;
	wire [31:0] mcycleh;
	wire [31:0] minstretl_ns;
	wire [31:0] minstretl;
	wire [31:0] minstreth_ns;
	wire [31:0] minstreth;
	wire [31:0] micect_ns;
	wire [31:0] micect;
	wire [31:0] miccmect_ns;
	wire [31:0] miccmect;
	wire [31:0] mdccmect_ns;
	wire [31:0] mdccmect;
	wire [26:0] micect_inc;
	wire [26:0] miccmect_inc;
	wire [26:0] mdccmect_inc;
	wire [31:0] mscratch;
	wire [31:0] mhpmc3;
	wire [31:0] mhpmc3_ns;
	wire [31:0] mhpmc4;
	wire [31:0] mhpmc4_ns;
	wire [31:0] mhpmc5;
	wire [31:0] mhpmc5_ns;
	wire [31:0] mhpmc6;
	wire [31:0] mhpmc6_ns;
	wire [31:0] mhpmc3h;
	wire [31:0] mhpmc3h_ns;
	wire [31:0] mhpmc4h;
	wire [31:0] mhpmc4h_ns;
	wire [31:0] mhpmc5h;
	wire [31:0] mhpmc5h_ns;
	wire [31:0] mhpmc6h;
	wire [31:0] mhpmc6h_ns;
	wire [9:0] mhpme3;
	wire [9:0] mhpme4;
	wire [9:0] mhpme5;
	wire [9:0] mhpme6;
	wire [31:0] mrac;
	wire [9:2] meihap;
	wire [31:10] meivt;
	wire [3:0] meicurpl_ns;
	wire [3:0] meicurpl;
	wire [3:0] meicidpl_ns;
	wire [3:0] meicidpl;
	wire [3:0] meipt_ns;
	wire [3:0] meipt;
	wire [31:0] mdseac;
	wire mdseac_locked_ns;
	wire mdseac_locked_f;
	wire mdseac_en;
	wire nmi_lsu_detected;
	wire [31:1] mepc_ns;
	wire [31:1] mepc;
	wire [31:1] dpc_ns;
	wire [31:1] dpc;
	wire [31:0] mcause_ns;
	wire [31:0] mcause;
	wire [3:0] mscause_ns;
	wire [3:0] mscause;
	wire [3:0] mscause_type;
	wire [31:0] mtval_ns;
	wire [31:0] mtval;
	wire dec_pause_state_f;
	wire dec_tlu_wr_pause_r_d1;
	wire pause_expired_r;
	wire pause_expired_wb;
	wire tlu_flush_lower_r;
	wire tlu_flush_lower_r_d1;
	wire [31:1] tlu_flush_path_r;
	wire [31:1] tlu_flush_path_r_d1;
	wire i0_valid_wb;
	wire tlu_i0_commit_cmt;
	wire [31:1] vectored_path;
	wire [31:1] interrupt_path;
	wire [16:0] dicawics_ns;
	wire [16:0] dicawics;
	wire wr_dicawics_r;
	wire wr_dicad0_r;
	wire wr_dicad1_r;
	wire wr_dicad0h_r;
	wire [31:0] dicad0_ns;
	wire [31:0] dicad0;
	wire [31:0] dicad0h_ns;
	wire [31:0] dicad0h;
	wire [6:0] dicad1_ns;
	wire [6:0] dicad1_raw;
	wire [31:0] dicad1;
	wire ebreak_r;
	wire ebreak_to_debug_mode_r;
	wire ecall_r;
	wire illegal_r;
	wire mret_r;
	wire inst_acc_r;
	wire fence_i_r;
	wire ic_perr_r;
	wire iccm_sbecc_r;
	wire ebreak_to_debug_mode_r_d1;
	wire kill_ebreak_count_r;
	wire inst_acc_second_r;
	wire ce_int_ready;
	wire ext_int_ready;
	wire timer_int_ready;
	wire soft_int_ready;
	wire int_timer0_int_ready;
	wire int_timer1_int_ready;
	wire mhwakeup_ready;
	wire take_ext_int;
	wire take_ce_int;
	wire take_timer_int;
	wire take_soft_int;
	wire take_int_timer0_int;
	wire take_int_timer1_int;
	wire take_nmi;
	wire take_nmi_r_d1;
	wire int_timer0_int_possible;
	wire int_timer1_int_possible;
	wire i0_exception_valid_r;
	wire interrupt_valid_r;
	wire i0_exception_valid_r_d1;
	wire interrupt_valid_r_d1;
	wire exc_or_int_valid_r;
	wire exc_or_int_valid_r_d1;
	wire mdccme_ce_req;
	wire miccme_ce_req;
	wire mice_ce_req;
	wire synchronous_flush_r;
	wire [4:0] exc_cause_r;
	wire [4:0] exc_cause_wb;
	wire mcyclel_cout;
	wire mcyclel_cout_f;
	wire mcyclela_cout;
	wire [31:0] mcyclel_inc;
	wire [31:0] mcycleh_inc;
	wire minstretl_cout;
	wire minstretl_cout_f;
	wire minstret_enable;
	wire minstretl_cout_ns;
	wire minstretl_couta;
	wire [31:0] minstretl_inc;
	wire [31:0] minstretl_read;
	wire [31:0] minstreth_inc;
	wire [31:0] minstreth_read;
	wire [31:1] pc_r;
	wire [31:1] pc_r_d1;
	wire [31:1] npc_r;
	wire [31:1] npc_r_d1;
	wire valid_csr;
	wire rfpc_i0_r;
	wire lsu_i0_rfnpc_r;
	wire dec_tlu_br0_error_r;
	wire dec_tlu_br0_start_error_r;
	wire dec_tlu_br0_v_r;
	wire lsu_i0_exc_r;
	wire lsu_i0_exc_r_raw;
	wire lsu_exc_ma_r;
	wire lsu_exc_acc_r;
	wire lsu_exc_st_r;
	wire lsu_exc_valid_r;
	wire lsu_exc_valid_r_raw;
	wire lsu_exc_valid_r_d1;
	wire lsu_i0_exc_r_d1;
	wire block_interrupts;
	wire i0_trigger_eval_r;
	wire request_debug_mode_r;
	wire request_debug_mode_r_d1;
	wire request_debug_mode_done;
	wire request_debug_mode_done_f;
	wire take_halt;
	wire halt_taken;
	wire halt_taken_f;
	wire internal_dbg_halt_mode;
	wire dbg_tlu_halted_f;
	wire take_reset;
	wire dbg_tlu_halted;
	wire core_empty;
	wire lsu_idle_any_f;
	wire ifu_miss_state_idle_f;
	wire resume_ack_ns;
	wire debug_halt_req_f;
	wire debug_resume_req_f_raw;
	wire debug_resume_req_f;
	wire enter_debug_halt_req;
	wire dcsr_single_step_done;
	wire dcsr_single_step_done_f;
	wire debug_halt_req_d1;
	wire debug_halt_req_ns;
	wire dcsr_single_step_running;
	wire dcsr_single_step_running_f;
	wire internal_dbg_halt_timers;
	wire [3:0] i0_trigger_r;
	wire [3:0] trigger_action;
	wire [3:0] trigger_enabled;
	wire [3:0] i0_trigger_chain_masked_r;
	wire i0_trigger_hit_r;
	wire i0_trigger_hit_raw_r;
	wire i0_trigger_action_r;
	wire trigger_hit_r_d1;
	wire mepc_trigger_hit_sel_pc_r;
	wire [3:0] update_hit_bit_r;
	wire [3:0] i0_iside_trigger_has_pri_r;
	wire [3:0] i0trigger_qual_r;
	wire [3:0] i0_lsu_trigger_has_pri_r;
	wire cpu_halt_status;
	wire cpu_halt_ack;
	wire cpu_run_ack;
	wire ext_halt_pulse;
	wire i_cpu_halt_req_d1;
	wire i_cpu_run_req_d1;
	wire inst_acc_r_raw;
	wire trigger_hit_dmode_r;
	wire trigger_hit_dmode_r_d1;
	wire [9:0] mcgc;
	wire [9:0] mcgc_ns;
	wire [9:0] mcgc_int;
	wire [18:0] mfdc;
	wire i_cpu_halt_req_sync_qual;
	wire i_cpu_run_req_sync_qual;
	wire pmu_fw_halt_req_ns;
	wire pmu_fw_halt_req_f;
	wire int_timer_stalled;
	wire fw_halt_req;
	wire enter_pmu_fw_halt_req;
	wire pmu_fw_tlu_halted;
	wire pmu_fw_tlu_halted_f;
	wire internal_pmu_fw_halt_mode;
	wire internal_pmu_fw_halt_mode_f;
	wire int_timer0_int_hold;
	wire int_timer1_int_hold;
	wire int_timer0_int_hold_f;
	wire int_timer1_int_hold_f;
	wire nmi_int_delayed;
	wire nmi_int_detected;
	wire [3:0] trigger_execute;
	wire [3:0] trigger_data;
	wire [3:0] trigger_store;
	wire dec_tlu_pmu_fw_halted;
	wire mpc_run_state_ns;
	wire debug_brkpt_status_ns;
	wire mpc_debug_halt_ack_ns;
	wire mpc_debug_run_ack_ns;
	wire dbg_halt_state_ns;
	wire dbg_run_state_ns;
	wire dbg_halt_state_f;
	wire mpc_debug_halt_req_sync_f;
	wire mpc_debug_run_req_sync_f;
	wire mpc_halt_state_f;
	wire mpc_halt_state_ns;
	wire mpc_run_state_f;
	wire debug_brkpt_status_f;
	wire mpc_debug_halt_ack_f;
	wire mpc_debug_run_ack_f;
	wire dbg_run_state_f;
	wire mpc_debug_halt_req_sync_pulse;
	wire mpc_debug_run_req_sync_pulse;
	wire debug_brkpt_valid;
	wire debug_halt_req;
	wire debug_resume_req;
	wire dec_tlu_mpc_halted_only_ns;
	wire take_ext_int_start;
	wire ext_int_freeze;
	wire take_ext_int_start_d1;
	wire take_ext_int_start_d2;
	wire take_ext_int_start_d3;
	wire ext_int_freeze_d1;
	wire csr_meicpct;
	wire ignore_ext_int_due_to_lsu_stall;
	wire mcause_sel_nmi_store;
	wire mcause_sel_nmi_load;
	wire mcause_sel_nmi_ext;
	wire fast_int_meicpct;
	wire [1:0] mcause_fir_error_type;
	wire dbg_halt_req_held_ns;
	wire dbg_halt_req_held;
	wire dbg_halt_req_final;
	wire iccm_repair_state_ns;
	wire iccm_repair_state_d1;
	wire iccm_repair_state_rfnpc;
	wire [31:0] dec_timer_rddata_d;
	wire dec_timer_read_d;
	wire dec_timer_t0_pulse;
	wire dec_timer_t1_pulse;
	wire csr_mitctl0;
	wire csr_mitctl1;
	wire csr_mitb0;
	wire csr_mitb1;
	wire csr_mitcnt0;
	wire csr_mitcnt1;
	wire nmi_int_sync;
	wire timer_int_sync;
	wire soft_int_sync;
	wire i_cpu_halt_req_sync;
	wire i_cpu_run_req_sync;
	wire mpc_debug_halt_req_sync;
	wire mpc_debug_run_req_sync;
	wire mpc_debug_halt_req_sync_raw;
	wire csr_wr_clk;
	wire e4e5_clk;
	wire e4_valid;
	wire e5_valid;
	wire e4e5_valid;
	wire internal_dbg_halt_mode_f;
	wire internal_dbg_halt_mode_f2;
	wire lsu_pmu_load_external_r;
	wire lsu_pmu_store_external_r;
	wire dec_tlu_flush_noredir_r_d1;
	wire dec_tlu_flush_pause_r_d1;
	wire lsu_single_ecc_error_r;
	wire [31:0] lsu_error_pkt_addr_r;
	wire mcyclel_cout_in;
	wire i0_valid_no_ebreak_ecall_r;
	wire minstret_enable_f;
	wire sel_exu_npc_r;
	wire sel_flush_npc_r;
	wire sel_hold_npc_r;
	wire pc0_valid_r;
	wire [15:0] mfdc_int;
	wire [15:0] mfdc_ns;
	wire [31:0] mrac_in;
	wire [31:27] csr_sat;
	wire [8:6] dcsr_cause;
	wire enter_debug_halt_req_le;
	wire dcsr_cause_upgradeable;
	wire icache_rd_valid;
	wire icache_wr_valid;
	wire icache_rd_valid_f;
	wire icache_wr_valid_f;
	wire [3:0] mhpmc_inc_r;
	wire [3:0] mhpmc_inc_r_d1;
	wire [39:0] mhpme_vec;
	wire mhpmc3_wr_en0;
	wire mhpmc3_wr_en1;
	wire mhpmc3_wr_en;
	wire mhpmc4_wr_en0;
	wire mhpmc4_wr_en1;
	wire mhpmc4_wr_en;
	wire mhpmc5_wr_en0;
	wire mhpmc5_wr_en1;
	wire mhpmc5_wr_en;
	wire mhpmc6_wr_en0;
	wire mhpmc6_wr_en1;
	wire mhpmc6_wr_en;
	wire mhpmc3h_wr_en0;
	wire mhpmc3h_wr_en;
	wire mhpmc4h_wr_en0;
	wire mhpmc4h_wr_en;
	wire mhpmc5h_wr_en0;
	wire mhpmc5h_wr_en;
	wire mhpmc6h_wr_en0;
	wire mhpmc6h_wr_en;
	wire [63:0] mhpmc3_incr;
	wire [63:0] mhpmc4_incr;
	wire [63:0] mhpmc5_incr;
	wire [63:0] mhpmc6_incr;
	wire perfcnt_halted_d1;
	wire zero_event_r;
	wire [3:0] perfcnt_during_sleep;
	wire [9:0] event_r;
	wire [3:0] pmu_i0_itype_qual;
	wire csr_mfdht;
	wire csr_mfdhs;
	wire csr_misa;
	wire csr_mvendorid;
	wire csr_marchid;
	wire csr_mimpid;
	wire csr_mhartid;
	wire csr_mstatus;
	wire csr_mtvec;
	wire csr_mip;
	wire csr_mie;
	wire csr_mcyclel;
	wire csr_mcycleh;
	wire csr_minstretl;
	wire csr_minstreth;
	wire csr_mscratch;
	wire csr_mepc;
	wire csr_mcause;
	wire csr_mscause;
	wire csr_mtval;
	wire csr_mrac;
	wire csr_dmst;
	wire csr_mdseac;
	wire csr_meihap;
	wire csr_meivt;
	wire csr_meipt;
	wire csr_meicurpl;
	wire csr_meicidpl;
	wire csr_dcsr;
	wire csr_mcgc;
	wire csr_mfdc;
	wire csr_dpc;
	wire csr_mtsel;
	wire csr_mtdata1;
	wire csr_mtdata2;
	wire csr_mhpmc3;
	wire csr_mhpmc4;
	wire csr_mhpmc5;
	wire csr_mhpmc6;
	wire csr_mhpmc3h;
	wire csr_mhpmc4h;
	wire csr_mhpmc5h;
	wire csr_mhpmc6h;
	wire csr_mhpme3;
	wire csr_mhpme4;
	wire csr_mhpme5;
	wire csr_mhpme6;
	wire csr_mcountinhibit;
	wire csr_mpmc;
	wire csr_micect;
	wire csr_miccmect;
	wire csr_mdccmect;
	wire csr_dicawics;
	wire csr_dicad0h;
	wire csr_dicad0;
	wire csr_dicad1;
	wire csr_dicago;
	wire presync;
	wire postsync;
	wire legal;
	wire dec_csr_wen_r_mod;
	wire flush_clkvalid;
	wire sel_fir_addr;
	wire wr_mie_r;
	wire mtval_capture_pc_r;
	wire mtval_capture_pc_plus2_r;
	wire mtval_capture_inst_r;
	wire mtval_capture_lsu_r;
	wire mtval_clear_r;
	wire wr_mcgc_r;
	wire wr_mfdc_r;
	wire wr_mdeau_r;
	wire trigger_hit_for_dscr_cause_r_d1;
	wire conditionally_illegal;
	wire [3:0] ifu_mscause;
	wire ifu_ic_error_start_f;
	wire ifu_iccm_rd_ecc_single_err_f;
	eb1_dec_timer_ctl #(.pt(pt)) int_timers(
		.clk(clk),
		.free_l2clk(free_l2clk),
		.csr_wr_clk(csr_wr_clk),
		.rst_l(rst_l),
		.dec_csr_wen_r_mod(dec_csr_wen_r_mod),
		.dec_csr_wraddr_r(dec_csr_wraddr_r),
		.dec_csr_wrdata_r(dec_csr_wrdata_r),
		.csr_mitctl0(csr_mitctl0),
		.csr_mitctl1(csr_mitctl1),
		.csr_mitb0(csr_mitb0),
		.csr_mitb1(csr_mitb1),
		.csr_mitcnt0(csr_mitcnt0),
		.csr_mitcnt1(csr_mitcnt1),
		.dec_pause_state(dec_pause_state),
		.dec_tlu_pmu_fw_halted(dec_tlu_pmu_fw_halted),
		.internal_dbg_halt_timers(internal_dbg_halt_timers),
		.dec_timer_rddata_d(dec_timer_rddata_d),
		.dec_timer_read_d(dec_timer_read_d),
		.dec_timer_t0_pulse(dec_timer_t0_pulse),
		.dec_timer_t1_pulse(dec_timer_t1_pulse),
		.scan_mode(scan_mode)
	);
	assign clk_override = dec_tlu_dec_clk_override;
	rvsyncss #(.WIDTH(7)) syncro_ff(
		.rst_l(rst_l),
		.clk(free_clk),
		.din({nmi_int, timer_int, soft_int, i_cpu_halt_req, i_cpu_run_req, mpc_debug_halt_req, mpc_debug_run_req}),
		.dout({nmi_int_sync, timer_int_sync, soft_int_sync, i_cpu_halt_req_sync, i_cpu_run_req_sync, mpc_debug_halt_req_sync_raw, mpc_debug_run_req_sync})
	);
	rvoclkhdr csrwr_r_cgc(
		.en(dec_csr_wen_r_mod | clk_override),
		.l1clk(csr_wr_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign e4_valid = dec_tlu_i0_valid_r;
	assign e4e5_valid = e4_valid | e5_valid;
	assign flush_clkvalid = ((((((((internal_dbg_halt_mode_f | i_cpu_run_req_d1) | interrupt_valid_r) | interrupt_valid_r_d1) | reset_delayed) | pause_expired_r) | pause_expired_wb) | ic_perr_r) | iccm_sbecc_r) | clk_override;
	rvoclkhdr e4e5_cgc(
		.en(e4e5_valid | clk_override),
		.l1clk(e4e5_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr e4e5_int_cgc(
		.en(e4e5_valid | flush_clkvalid),
		.l1clk(e4e5_int_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvdffie #(.WIDTH(11)) freeff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({ifu_ic_error_start, ifu_iccm_rd_ecc_single_err, iccm_repair_state_ns, e4_valid, internal_dbg_halt_mode, lsu_pmu_load_external_m, lsu_pmu_store_external_m, tlu_flush_lower_r, tlu_i0_kill_writeb_r, internal_dbg_halt_mode_f, force_halt}),
		.dout({ifu_ic_error_start_f, ifu_iccm_rd_ecc_single_err_f, iccm_repair_state_d1, e5_valid, internal_dbg_halt_mode_f, lsu_pmu_load_external_r, lsu_pmu_store_external_r, tlu_flush_lower_r_d1, dec_tlu_i0_kill_writeb_wb, internal_dbg_halt_mode_f2, dec_tlu_force_halt})
	);
	assign dec_tlu_i0_kill_writeb_r = tlu_i0_kill_writeb_r;
	assign nmi_int_detected = (((nmi_int_sync & ~nmi_int_delayed) | nmi_lsu_detected) | (nmi_int_detected_f & ~take_nmi_r_d1)) | nmi_fir_type;
	assign nmi_lsu_load_type = ((nmi_lsu_detected & lsu_imprecise_error_load_any) & ~(nmi_int_detected_f & ~take_nmi_r_d1)) | (nmi_lsu_load_type_f & ~take_nmi_r_d1);
	assign nmi_lsu_store_type = ((nmi_lsu_detected & lsu_imprecise_error_store_any) & ~(nmi_int_detected_f & ~take_nmi_r_d1)) | (nmi_lsu_store_type_f & ~take_nmi_r_d1);
	assign nmi_fir_type = (~nmi_int_detected_f & take_ext_int_start_d3) & |lsu_fir_error[1:0];
	assign nmi_lsu_detected = (~mdseac_locked_f & (lsu_imprecise_error_load_any | lsu_imprecise_error_store_any)) & ~nmi_fir_type;
	localparam MSTATUS_MIE = 0;
	localparam MIP_MCEIP = 5;
	localparam MIP_MITIP0 = 4;
	localparam MIP_MITIP1 = 3;
	localparam MIP_MEIP = 2;
	localparam MIP_MTIP = 1;
	localparam MIP_MSIP = 0;
	localparam MIE_MCEIE = 5;
	localparam MIE_MITIE0 = 4;
	localparam MIE_MITIE1 = 3;
	localparam MIE_MEIE = 2;
	localparam MIE_MTIE = 1;
	localparam MIE_MSIE = 0;
	localparam DCSR_EBREAKM = 15;
	localparam DCSR_STEPIE = 11;
	localparam DCSR_STOPC = 10;
	localparam DCSR_STEP = 2;
	assign reset_delayed = reset_detect ^ reset_detected;
	assign mpc_debug_halt_req_sync = mpc_debug_halt_req_sync_raw & ~ext_int_freeze_d1;
	rvdffie #(.WIDTH(16)) mpvhalt_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({1'b1, reset_detect, nmi_int_sync, nmi_int_detected, nmi_lsu_load_type, nmi_lsu_store_type, mpc_debug_halt_req_sync, mpc_debug_run_req_sync, mpc_halt_state_ns, mpc_run_state_ns, debug_brkpt_status_ns, mpc_debug_halt_ack_ns, mpc_debug_run_ack_ns, dbg_halt_state_ns, dbg_run_state_ns, dec_tlu_mpc_halted_only_ns}),
		.dout({reset_detect, reset_detected, nmi_int_delayed, nmi_int_detected_f, nmi_lsu_load_type_f, nmi_lsu_store_type_f, mpc_debug_halt_req_sync_f, mpc_debug_run_req_sync_f, mpc_halt_state_f, mpc_run_state_f, debug_brkpt_status_f, mpc_debug_halt_ack_f, mpc_debug_run_ack_f, dbg_halt_state_f, dbg_run_state_f, dec_tlu_mpc_halted_only})
	);
	assign mpc_debug_halt_req_sync_pulse = mpc_debug_halt_req_sync & ~mpc_debug_halt_req_sync_f;
	assign mpc_debug_run_req_sync_pulse = mpc_debug_run_req_sync & ~mpc_debug_run_req_sync_f;
	assign mpc_halt_state_ns = ((mpc_halt_state_f | mpc_debug_halt_req_sync_pulse) | (reset_delayed & ~mpc_reset_run_req)) & ~mpc_debug_run_req_sync;
	assign mpc_run_state_ns = (mpc_run_state_f | (mpc_debug_run_req_sync_pulse & ~mpc_debug_run_ack_f)) & (internal_dbg_halt_mode_f & ~dcsr_single_step_running_f);
	assign dbg_halt_state_ns = (dbg_halt_state_f | (((dbg_halt_req_final | dcsr_single_step_done_f) | trigger_hit_dmode_r_d1) | ebreak_to_debug_mode_r_d1)) & ~dbg_resume_req;
	assign dbg_run_state_ns = (dbg_run_state_f | dbg_resume_req) & (internal_dbg_halt_mode_f & ~dcsr_single_step_running_f);
	assign dec_tlu_mpc_halted_only_ns = ~dbg_halt_state_f & mpc_halt_state_f;
	assign debug_brkpt_valid = ebreak_to_debug_mode_r_d1 | trigger_hit_dmode_r_d1;
	assign debug_brkpt_status_ns = (debug_brkpt_valid | debug_brkpt_status_f) & (internal_dbg_halt_mode & ~dcsr_single_step_running_f);
	assign mpc_debug_halt_ack_ns = ((mpc_halt_state_f & internal_dbg_halt_mode_f) & mpc_debug_halt_req_sync) & core_empty;
	assign mpc_debug_run_ack_ns = ((mpc_debug_run_req_sync & ~dbg_halt_state_ns) & ~mpc_debug_halt_req_sync) | (mpc_debug_run_ack_f & mpc_debug_run_req_sync);
	assign mpc_debug_halt_ack = mpc_debug_halt_ack_f;
	assign mpc_debug_run_ack = mpc_debug_run_ack_f;
	assign debug_brkpt_status = debug_brkpt_status_f;
	assign dbg_halt_req_held_ns = (dbg_halt_req | dbg_halt_req_held) & ext_int_freeze_d1;
	assign dbg_halt_req_final = (dbg_halt_req | dbg_halt_req_held) & ~ext_int_freeze_d1;
	assign debug_halt_req = (((dbg_halt_req_final | mpc_debug_halt_req_sync) | (reset_delayed & ~mpc_reset_run_req)) & ~internal_dbg_halt_mode_f) & ~ext_int_freeze_d1;
	assign debug_resume_req = ~debug_resume_req_f & ((mpc_run_state_ns & ~dbg_halt_state_ns) | (dbg_run_state_ns & ~mpc_halt_state_ns));
	assign take_halt = (((((debug_halt_req_f | pmu_fw_halt_req_f) & ~synchronous_flush_r) & ~mret_r) & ~halt_taken_f) & ~dec_tlu_flush_noredir_r_d1) & ~take_reset;
	assign halt_taken = ((dec_tlu_flush_noredir_r_d1 & ~dec_tlu_flush_pause_r_d1) & ~take_ext_int_start_d1) | (((halt_taken_f & ~dbg_tlu_halted_f) & ~pmu_fw_tlu_halted_f) & ~interrupt_valid_r_d1);
	assign core_empty = force_halt | ((((((lsu_idle_any & lsu_idle_any_f) & ifu_miss_state_idle) & ifu_miss_state_idle_f) & ~debug_halt_req) & ~debug_halt_req_d1) & ~dec_div_active);
	assign dec_tlu_core_empty = core_empty;
	assign enter_debug_halt_req = (((~internal_dbg_halt_mode_f & debug_halt_req) | dcsr_single_step_done_f) | trigger_hit_dmode_r_d1) | ebreak_to_debug_mode_r_d1;
	assign internal_dbg_halt_mode = debug_halt_req_ns | (internal_dbg_halt_mode_f & ~(debug_resume_req_f & ~dcsr[DCSR_STEP]));
	assign allow_dbg_halt_csr_write = internal_dbg_halt_mode_f & ~dcsr_single_step_running_f;
	assign debug_halt_req_ns = enter_debug_halt_req | (debug_halt_req_f & ~dbg_tlu_halted);
	assign dbg_tlu_halted = ((debug_halt_req_f & core_empty) & halt_taken) | (dbg_tlu_halted_f & ~debug_resume_req_f);
	assign resume_ack_ns = (debug_resume_req_f & dbg_tlu_halted_f) & dbg_run_state_ns;
	assign dcsr_single_step_done = ((dec_tlu_i0_valid_r & ~dec_tlu_dbg_halted) & dcsr[DCSR_STEP]) & ~rfpc_i0_r;
	assign dcsr_single_step_running = (debug_resume_req_f & dcsr[DCSR_STEP]) | (dcsr_single_step_running_f & ~dcsr_single_step_done_f);
	assign dbg_cmd_done_ns = dec_tlu_i0_valid_r & dec_tlu_dbg_halted;
	assign request_debug_mode_r = (trigger_hit_dmode_r | ebreak_to_debug_mode_r) | (request_debug_mode_r_d1 & ~dec_tlu_flush_lower_wb);
	assign request_debug_mode_done = (request_debug_mode_r_d1 | request_debug_mode_done_f) & ~dbg_tlu_halted_f;
	rvdffie #(.WIDTH(18)) halt_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({dec_tlu_flush_noredir_r, halt_taken, lsu_idle_any, ifu_miss_state_idle, dbg_tlu_halted, resume_ack_ns, debug_halt_req_ns, debug_resume_req, trigger_hit_dmode_r, dcsr_single_step_done, debug_halt_req, dec_tlu_wr_pause_r, dec_pause_state, request_debug_mode_r, request_debug_mode_done, dcsr_single_step_running, dec_tlu_flush_pause_r, dbg_halt_req_held_ns}),
		.dout({dec_tlu_flush_noredir_r_d1, halt_taken_f, lsu_idle_any_f, ifu_miss_state_idle_f, dbg_tlu_halted_f, dec_tlu_resume_ack, debug_halt_req_f, debug_resume_req_f_raw, trigger_hit_dmode_r_d1, dcsr_single_step_done_f, debug_halt_req_d1, dec_tlu_wr_pause_r_d1, dec_pause_state_f, request_debug_mode_r_d1, request_debug_mode_done_f, dcsr_single_step_running_f, dec_tlu_flush_pause_r_d1, dbg_halt_req_held})
	);
	assign debug_resume_req_f = debug_resume_req_f_raw & ~dbg_halt_req;
	assign dec_tlu_debug_stall = debug_halt_req_f;
	assign dec_tlu_dbg_halted = dbg_tlu_halted_f;
	assign dec_tlu_debug_mode = internal_dbg_halt_mode_f;
	assign dec_tlu_pmu_fw_halted = pmu_fw_tlu_halted_f;
	assign dec_tlu_flush_noredir_r = (((take_halt | (fence_i_r & internal_dbg_halt_mode)) | dec_tlu_flush_pause_r) | (i0_trigger_hit_r & trigger_hit_dmode_r)) | take_ext_int_start;
	assign dec_tlu_flush_extint = take_ext_int_start;
	assign dec_tlu_flush_pause_r = (dec_tlu_wr_pause_r_d1 & ~interrupt_valid_r) & ~take_ext_int_start;
	assign pause_expired_r = (((((~dec_pause_state & dec_pause_state_f) & ~(((((((ext_int_ready | ce_int_ready) | timer_int_ready) | soft_int_ready) | int_timer0_int_hold_f) | int_timer1_int_hold_f) | nmi_int_detected) | ext_int_freeze_d1)) & ~interrupt_valid_r_d1) & ~debug_halt_req_f) & ~pmu_fw_halt_req_f) & ~halt_taken_f;
	assign dec_tlu_flush_leak_one_r = ((dec_tlu_flush_lower_r & dcsr[DCSR_STEP]) & (dec_tlu_resume_ack | dcsr_single_step_running)) & ~dec_tlu_flush_noredir_r;
	assign dec_tlu_flush_err_r = dec_tlu_flush_lower_r & (ic_perr_r | iccm_sbecc_r);
	assign dec_dbg_cmd_done = dbg_cmd_done_ns;
	assign dec_dbg_cmd_fail = illegal_r & dec_dbg_cmd_done;
	localparam MTDATA1_DMODE = 9;
	localparam MTDATA1_SEL = 7;
	localparam MTDATA1_ACTION = 6;
	localparam MTDATA1_CHAIN = 5;
	localparam MTDATA1_MATCH = 4;
	localparam MTDATA1_M_ENABLED = 3;
	localparam MTDATA1_EXE = 2;
	localparam MTDATA1_ST = 1;
	localparam MTDATA1_LD = 0;
	assign trigger_execute[3:0] = {mtdata1_t3[MTDATA1_EXE], mtdata1_t2[MTDATA1_EXE], mtdata1_t1[MTDATA1_EXE], mtdata1_t0[MTDATA1_EXE]};
	assign trigger_data[3:0] = {mtdata1_t3[MTDATA1_SEL], mtdata1_t2[MTDATA1_SEL], mtdata1_t1[MTDATA1_SEL], mtdata1_t0[MTDATA1_SEL]};
	assign trigger_store[3:0] = {mtdata1_t3[MTDATA1_ST], mtdata1_t2[MTDATA1_ST], mtdata1_t1[MTDATA1_ST], mtdata1_t0[MTDATA1_ST]};
	assign trigger_enabled[3:0] = {(mtdata1_t3[MTDATA1_ACTION] | mstatus[MSTATUS_MIE]) & mtdata1_t3[MTDATA1_M_ENABLED], (mtdata1_t2[MTDATA1_ACTION] | mstatus[MSTATUS_MIE]) & mtdata1_t2[MTDATA1_M_ENABLED], (mtdata1_t1[MTDATA1_ACTION] | mstatus[MSTATUS_MIE]) & mtdata1_t1[MTDATA1_M_ENABLED], (mtdata1_t0[MTDATA1_ACTION] | mstatus[MSTATUS_MIE]) & mtdata1_t0[MTDATA1_M_ENABLED]};
	assign i0_iside_trigger_has_pri_r[3:0] = ~(((trigger_execute[3:0] & trigger_data[3:0]) & {4 {inst_acc_r_raw}}) | {4 {exu_i0_br_error_r | exu_i0_br_start_error_r}});
	assign i0_lsu_trigger_has_pri_r[3:0] = ~((trigger_store[3:0] & trigger_data[3:0]) & {4 {lsu_i0_exc_r_raw}});
	assign i0_trigger_eval_r = dec_tlu_i0_valid_r;
	assign i0trigger_qual_r[3:0] = ((({4 {i0_trigger_eval_r}} & dec_tlu_packet_r[11:8]) & i0_iside_trigger_has_pri_r[3:0]) & i0_lsu_trigger_has_pri_r[3:0]) & trigger_enabled[3:0];
	assign i0_trigger_r[3:0] = ~{4 {dec_tlu_flush_lower_wb | dec_tlu_dbg_halted}} & i0trigger_qual_r[3:0];
	assign i0_trigger_chain_masked_r[3:0] = {i0_trigger_r[3] & (~mtdata1_t2[MTDATA1_CHAIN] | i0_trigger_r[2]), i0_trigger_r[2] & (~mtdata1_t2[MTDATA1_CHAIN] | i0_trigger_r[3]), i0_trigger_r[1] & (~mtdata1_t0[MTDATA1_CHAIN] | i0_trigger_r[0]), i0_trigger_r[0] & (~mtdata1_t0[MTDATA1_CHAIN] | i0_trigger_r[1])};
	assign i0_trigger_hit_raw_r = |i0_trigger_chain_masked_r[3:0];
	assign i0_trigger_hit_r = i0_trigger_hit_raw_r;
	assign trigger_action[3:0] = {mtdata1_t3[MTDATA1_ACTION] & mtdata1_t3[MTDATA1_DMODE], (mtdata1_t2[MTDATA1_ACTION] & mtdata1_t2[MTDATA1_DMODE]) & ~mtdata1_t2[MTDATA1_CHAIN], mtdata1_t1[MTDATA1_ACTION] & mtdata1_t1[MTDATA1_DMODE], (mtdata1_t0[MTDATA1_ACTION] & mtdata1_t0[MTDATA1_DMODE]) & ~mtdata1_t0[MTDATA1_CHAIN]};
	assign update_hit_bit_r[3:0] = {4 {|i0_trigger_r[3:0] & ~rfpc_i0_r}} & {i0_trigger_chain_masked_r[3], i0_trigger_r[2], i0_trigger_chain_masked_r[1], i0_trigger_r[0]};
	assign i0_trigger_action_r = |(i0_trigger_chain_masked_r[3:0] & trigger_action[3:0]);
	assign trigger_hit_dmode_r = i0_trigger_hit_r & i0_trigger_action_r;
	assign mepc_trigger_hit_sel_pc_r = i0_trigger_hit_r & ~trigger_hit_dmode_r;
	assign i_cpu_halt_req_sync_qual = (i_cpu_halt_req_sync & ~dec_tlu_debug_mode) & ~ext_int_freeze_d1;
	assign i_cpu_run_req_sync_qual = ((i_cpu_run_req_sync & ~dec_tlu_debug_mode) & pmu_fw_tlu_halted_f) & ~ext_int_freeze_d1;
	rvdffie #(.WIDTH(10)) exthaltff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({i_cpu_halt_req_sync_qual, i_cpu_run_req_sync_qual, cpu_halt_status, cpu_halt_ack, cpu_run_ack, internal_pmu_fw_halt_mode, pmu_fw_halt_req_ns, pmu_fw_tlu_halted, int_timer0_int_hold, int_timer1_int_hold}),
		.dout({i_cpu_halt_req_d1, i_cpu_run_req_d1_raw, o_cpu_halt_status, o_cpu_halt_ack, o_cpu_run_ack, internal_pmu_fw_halt_mode_f, pmu_fw_halt_req_f, pmu_fw_tlu_halted_f, int_timer0_int_hold_f, int_timer1_int_hold_f})
	);
	assign ext_halt_pulse = i_cpu_halt_req_sync_qual & ~i_cpu_halt_req_d1;
	assign enter_pmu_fw_halt_req = ext_halt_pulse | fw_halt_req;
	assign pmu_fw_halt_req_ns = (enter_pmu_fw_halt_req | (pmu_fw_halt_req_f & ~pmu_fw_tlu_halted)) & ~debug_halt_req_f;
	assign internal_pmu_fw_halt_mode = pmu_fw_halt_req_ns | ((internal_pmu_fw_halt_mode_f & ~i_cpu_run_req_d1) & ~debug_halt_req_f);
	assign pmu_fw_tlu_halted = ((((pmu_fw_halt_req_f & core_empty) & halt_taken) & ~enter_debug_halt_req) | (pmu_fw_tlu_halted_f & ~i_cpu_run_req_d1)) & ~debug_halt_req_f;
	assign cpu_halt_ack = (i_cpu_halt_req_d1 & pmu_fw_tlu_halted_f) | (o_cpu_halt_ack & i_cpu_halt_req_sync);
	assign cpu_halt_status = (pmu_fw_tlu_halted_f & ~i_cpu_run_req_d1) | ((o_cpu_halt_status & ~i_cpu_run_req_d1) & ~internal_dbg_halt_mode_f);
	assign cpu_run_ack = ((~pmu_fw_tlu_halted_f & i_cpu_run_req_sync) | (o_cpu_halt_status & i_cpu_run_req_d1_raw)) | (o_cpu_run_ack & i_cpu_run_req_sync);
	assign debug_mode_status = internal_dbg_halt_mode_f;
	assign o_debug_mode_status = debug_mode_status;
	assign i_cpu_run_req_d1 = i_cpu_run_req_d1_raw | (((((((nmi_int_detected | timer_int_ready) | soft_int_ready) | int_timer0_int_hold_f) | int_timer1_int_hold_f) | (mhwakeup & mhwakeup_ready)) & o_cpu_halt_status) & ~i_cpu_halt_req_d1);
	assign lsu_single_ecc_error_r = lsu_single_ecc_error_incr;
	assign lsu_error_pkt_addr_r[31:0] = lsu_error_pkt_r[33:2];
	assign lsu_exc_valid_r_raw = lsu_error_pkt_r[0] & ~dec_tlu_flush_lower_wb;
	assign lsu_i0_exc_r_raw = lsu_error_pkt_r[0];
	assign lsu_i0_exc_r = ((lsu_i0_exc_r_raw & lsu_exc_valid_r_raw) & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	assign lsu_exc_valid_r = lsu_i0_exc_r;
	assign lsu_exc_ma_r = lsu_i0_exc_r & ~lsu_error_pkt_r[38];
	assign lsu_exc_acc_r = lsu_i0_exc_r & lsu_error_pkt_r[38];
	assign lsu_exc_st_r = lsu_i0_exc_r & lsu_error_pkt_r[39];
	assign lsu_i0_rfnpc_r = (dec_tlu_i0_valid_r & ~i0_trigger_hit_r) & (~lsu_error_pkt_r[39] & lsu_error_pkt_r[1]);
	assign tlu_i0_commit_cmt = (((((dec_tlu_i0_valid_r & ~rfpc_i0_r) & ~lsu_i0_exc_r) & ~inst_acc_r) & ~dec_tlu_dbg_halted) & ~request_debug_mode_r_d1) & ~i0_trigger_hit_r;
	assign tlu_i0_kill_writeb_r = (((rfpc_i0_r | lsu_i0_exc_r) | inst_acc_r) | (illegal_r & dec_tlu_dbg_halted)) | i0_trigger_hit_r;
	assign dec_tlu_i0_commit_cmt = tlu_i0_commit_cmt;
	assign rfpc_i0_r = ((((dec_tlu_i0_valid_r & ~tlu_flush_lower_r_d1) & (exu_i0_br_error_r | exu_i0_br_start_error_r)) | ((ic_perr_r | iccm_sbecc_r) & ~ext_int_freeze_d1)) & ~i0_trigger_hit_r) & ~lsu_i0_rfnpc_r;
	assign iccm_repair_state_ns = iccm_sbecc_r | (iccm_repair_state_d1 & ~dec_tlu_flush_lower_r);
	localparam MCPC = 12'h7c2;
	assign iccm_repair_state_rfnpc = (tlu_i0_commit_cmt & iccm_repair_state_d1) & ~(((((ebreak_r | ecall_r) | mret_r) | take_reset) | illegal_r) | (dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCPC)));
	generate
		if (pt[2130-:5] == 1) begin
			assign dec_tlu_br0_error_r = (exu_i0_br_error_r & dec_tlu_i0_valid_r) & ~tlu_flush_lower_r_d1;
			assign dec_tlu_br0_start_error_r = (exu_i0_br_start_error_r & dec_tlu_i0_valid_r) & ~tlu_flush_lower_r_d1;
			assign dec_tlu_br0_v_r = ((exu_i0_br_valid_r & dec_tlu_i0_valid_r) & ~tlu_flush_lower_r_d1) & (~exu_i0_br_mp_r | ~exu_pmu_i0_br_ataken);
			assign dec_tlu_br0_r_pkt[5:4] = exu_i0_br_hist_r[1:0];
			assign dec_tlu_br0_r_pkt[3] = dec_tlu_br0_error_r;
			assign dec_tlu_br0_r_pkt[2] = dec_tlu_br0_start_error_r;
			assign dec_tlu_br0_r_pkt[6] = dec_tlu_br0_v_r;
			assign dec_tlu_br0_r_pkt[1] = exu_i0_br_way_r;
			assign dec_tlu_br0_r_pkt[0] = exu_i0_br_middle_r;
		end
		else begin
			assign dec_tlu_br0_error_r = 1'b0;
			assign dec_tlu_br0_start_error_r = 1'b0;
			assign dec_tlu_br0_v_r = 1'b0;
			assign dec_tlu_br0_r_pkt = {7 {1'sb0}};
		end
	endgenerate
	localparam [3:0] eb1_pkg_EBREAK = 4'b1000;
	assign ebreak_r = ((((dec_tlu_packet_r[3-:4] == eb1_pkg_EBREAK) & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & ~dcsr[DCSR_EBREAKM]) & ~rfpc_i0_r;
	localparam [3:0] eb1_pkg_ECALL = 4'b1001;
	assign ecall_r = (((dec_tlu_packet_r[3-:4] == eb1_pkg_ECALL) & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	assign illegal_r = ((~dec_tlu_packet_r[5] & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	localparam [3:0] eb1_pkg_MRET = 4'b1100;
	assign mret_r = (((dec_tlu_packet_r[3-:4] == eb1_pkg_MRET) & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	assign fence_i_r = ((dec_tlu_packet_r[12] & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	assign ic_perr_r = ((ifu_ic_error_start_f & ~ext_int_freeze_d1) & (~internal_dbg_halt_mode_f | dcsr_single_step_running)) & ~internal_pmu_fw_halt_mode_f;
	assign iccm_sbecc_r = ((ifu_iccm_rd_ecc_single_err_f & ~ext_int_freeze_d1) & (~internal_dbg_halt_mode_f | dcsr_single_step_running)) & ~internal_pmu_fw_halt_mode_f;
	assign inst_acc_r_raw = dec_tlu_packet_r[16] & dec_tlu_i0_valid_r;
	assign inst_acc_r = (inst_acc_r_raw & ~rfpc_i0_r) & ~i0_trigger_hit_r;
	assign inst_acc_second_r = dec_tlu_packet_r[15];
	assign ebreak_to_debug_mode_r = ((((dec_tlu_packet_r[3-:4] == eb1_pkg_EBREAK) & dec_tlu_i0_valid_r) & ~i0_trigger_hit_r) & dcsr[DCSR_EBREAKM]) & ~rfpc_i0_r;
	rvdff #(.WIDTH(1)) exctype_wb_ff(
		.rst_l(rst_l),
		.clk(e4e5_clk),
		.din(ebreak_to_debug_mode_r),
		.dout(ebreak_to_debug_mode_r_d1)
	);
	assign dec_tlu_fence_i_r = fence_i_r;
	assign i0_exception_valid_r = ((((ebreak_r | ecall_r) | illegal_r) | inst_acc_r) & ~rfpc_i0_r) & ~dec_tlu_dbg_halted;
	assign exc_cause_r[4:0] = (((((((((((((({5 {take_ext_int}} & 5'h0b) | ({5 {take_timer_int}} & 5'h07)) | ({5 {take_soft_int}} & 5'h03)) | ({5 {take_int_timer0_int}} & 5'h1d)) | ({5 {take_int_timer1_int}} & 5'h1c)) | ({5 {take_ce_int}} & 5'h1e)) | ({5 {illegal_r}} & 5'h02)) | ({5 {ecall_r}} & 5'h0b)) | ({5 {inst_acc_r}} & 5'h01)) | ({5 {ebreak_r | i0_trigger_hit_r}} & 5'h03)) | ({5 {lsu_exc_ma_r & ~lsu_exc_st_r}} & 5'h04)) | ({5 {lsu_exc_acc_r & ~lsu_exc_st_r}} & 5'h05)) | ({5 {lsu_exc_ma_r & lsu_exc_st_r}} & 5'h06)) | ({5 {lsu_exc_acc_r & lsu_exc_st_r}} & 5'h07)) & ~{5 {take_nmi}};
	assign mhwakeup_ready = ((~dec_csr_stall_int_ff & mstatus_mie_ns) & mip[MIP_MEIP]) & mie_ns[MIE_MEIE];
	assign ext_int_ready = (((~dec_csr_stall_int_ff & mstatus_mie_ns) & mip[MIP_MEIP]) & mie_ns[MIE_MEIE]) & ~ignore_ext_int_due_to_lsu_stall;
	assign ce_int_ready = ((~dec_csr_stall_int_ff & mstatus_mie_ns) & mip[MIP_MCEIP]) & mie_ns[MIE_MCEIE];
	assign soft_int_ready = ((~dec_csr_stall_int_ff & mstatus_mie_ns) & mip[MIP_MSIP]) & mie_ns[MIE_MSIE];
	assign timer_int_ready = ((~dec_csr_stall_int_ff & mstatus_mie_ns) & mip[MIP_MTIP]) & mie_ns[MIE_MTIE];
	assign int_timer0_int_possible = mstatus_mie_ns & mie_ns[MIE_MITIE0];
	assign int_timer0_int_ready = mip[MIP_MITIP0] & int_timer0_int_possible;
	assign int_timer1_int_possible = mstatus_mie_ns & mie_ns[MIE_MITIE1];
	assign int_timer1_int_ready = mip[MIP_MITIP1] & int_timer1_int_possible;
	assign int_timer_stalled = ((dec_csr_stall_int_ff | synchronous_flush_r) | exc_or_int_valid_r_d1) | mret_r;
	assign int_timer0_int_hold = (int_timer0_int_ready & (pmu_fw_tlu_halted_f | int_timer_stalled)) | ((((int_timer0_int_possible & int_timer0_int_hold_f) & ~interrupt_valid_r) & ~take_ext_int_start) & ~internal_dbg_halt_mode_f);
	assign int_timer1_int_hold = (int_timer1_int_ready & (pmu_fw_tlu_halted_f | int_timer_stalled)) | ((((int_timer1_int_possible & int_timer1_int_hold_f) & ~interrupt_valid_r) & ~take_ext_int_start) & ~internal_dbg_halt_mode_f);
	assign internal_dbg_halt_timers = internal_dbg_halt_mode_f & ~dcsr_single_step_running;
	assign block_interrupts = ((((((((internal_dbg_halt_mode & (~dcsr_single_step_running | dec_tlu_i0_valid_r)) | internal_pmu_fw_halt_mode) | i_cpu_halt_req_d1) | take_nmi) | ebreak_to_debug_mode_r) | synchronous_flush_r) | exc_or_int_valid_r_d1) | mret_r) | ext_int_freeze_d1;
	generate
		if (pt[1227-:5]) begin
			assign take_ext_int_start = ext_int_ready & ~block_interrupts;
			assign ext_int_freeze = ((take_ext_int_start | take_ext_int_start_d1) | take_ext_int_start_d2) | take_ext_int_start_d3;
			assign take_ext_int = take_ext_int_start_d3 & ~|lsu_fir_error[1:0];
			assign fast_int_meicpct = csr_meicpct & dec_csr_any_unq_d;
			assign ignore_ext_int_due_to_lsu_stall = lsu_fastint_stall_any;
		end
		else begin
			assign take_ext_int_start = 1'b0;
			assign ext_int_freeze = 1'b0;
			assign ext_int_freeze_d1 = 1'b0;
			assign take_ext_int_start_d1 = 1'b0;
			assign take_ext_int_start_d2 = 1'b0;
			assign take_ext_int_start_d3 = 1'b0;
			assign fast_int_meicpct = 1'b0;
			assign ignore_ext_int_due_to_lsu_stall = 1'b0;
			assign take_ext_int = ext_int_ready & ~block_interrupts;
		end
	endgenerate
	assign take_ce_int = (ce_int_ready & ~ext_int_ready) & ~block_interrupts;
	assign take_soft_int = ((soft_int_ready & ~ext_int_ready) & ~ce_int_ready) & ~block_interrupts;
	assign take_timer_int = (((timer_int_ready & ~soft_int_ready) & ~ext_int_ready) & ~ce_int_ready) & ~block_interrupts;
	assign take_int_timer0_int = (((((((int_timer0_int_ready | int_timer0_int_hold_f) & int_timer0_int_possible) & ~dec_csr_stall_int_ff) & ~timer_int_ready) & ~soft_int_ready) & ~ext_int_ready) & ~ce_int_ready) & ~block_interrupts;
	assign take_int_timer1_int = ((((((((int_timer1_int_ready | int_timer1_int_hold_f) & int_timer1_int_possible) & ~dec_csr_stall_int_ff) & ~(int_timer0_int_ready | int_timer0_int_hold_f)) & ~timer_int_ready) & ~soft_int_ready) & ~ext_int_ready) & ~ce_int_ready) & ~block_interrupts;
	assign take_reset = reset_delayed & mpc_reset_run_req;
	assign take_nmi = ((((((nmi_int_detected & ~internal_pmu_fw_halt_mode) & (~internal_dbg_halt_mode | (((dcsr_single_step_running_f & dcsr[DCSR_STEPIE]) & ~dec_tlu_i0_valid_r) & ~dcsr_single_step_done_f))) & ~synchronous_flush_r) & ~mret_r) & ~take_reset) & ~ebreak_to_debug_mode_r) & (~ext_int_freeze_d1 | (take_ext_int_start_d3 & |lsu_fir_error[1:0]));
	assign interrupt_valid_r = (((((take_ext_int | take_timer_int) | take_soft_int) | take_nmi) | take_ce_int) | take_int_timer0_int) | take_int_timer1_int;
	assign vectored_path[31:1] = {mtvec[30:1], 1'b0} + {25'b0000000000000000000000000, exc_cause_r[4:0], 1'b0};
	assign interrupt_path[31:1] = (take_nmi ? nmi_vec[31:1] : (mtvec[0] == 1'b1 ? vectored_path[31:1] : {mtvec[30:1], 1'b0}));
	assign sel_npc_r = (((lsu_i0_rfnpc_r | fence_i_r) | iccm_repair_state_rfnpc) | (i_cpu_run_req_d1 & ~interrupt_valid_r)) | (rfpc_i0_r & ~dec_tlu_i0_valid_r);
	assign sel_npc_resume = (i_cpu_run_req_d1 & pmu_fw_tlu_halted_f) | pause_expired_r;
	assign sel_fir_addr = take_ext_int_start_d3 & ~|lsu_fir_error[1:0];
	assign synchronous_flush_r = ((((((((i0_exception_valid_r | rfpc_i0_r) | lsu_exc_valid_r) | fence_i_r) | lsu_i0_rfnpc_r) | iccm_repair_state_rfnpc) | debug_resume_req_f) | sel_npc_resume) | dec_tlu_wr_pause_r_d1) | i0_trigger_hit_r;
	assign tlu_flush_lower_r = ((((interrupt_valid_r | mret_r) | synchronous_flush_r) | take_halt) | take_reset) | take_ext_int_start;
	assign tlu_flush_path_r[31:1] = (take_reset ? rst_vec[31:1] : ((((((({31 {sel_fir_addr}} & lsu_fir_addr[31:1]) | ({31 {~take_nmi & sel_npc_r}} & npc_r[31:1])) | ({31 {((~take_nmi & rfpc_i0_r) & dec_tlu_i0_valid_r) & ~sel_npc_r}} & dec_tlu_i0_pc_r[31:1])) | ({31 {interrupt_valid_r & ~sel_fir_addr}} & interrupt_path[31:1])) | ({31 {(((i0_exception_valid_r | lsu_exc_valid_r) | (i0_trigger_hit_r & ~trigger_hit_dmode_r)) & ~interrupt_valid_r) & ~sel_fir_addr}} & {mtvec[30:1], 1'b0})) | ({31 {~take_nmi & mret_r}} & mepc[31:1])) | ({31 {~take_nmi & debug_resume_req_f}} & dpc[31:1])) | ({31 {~take_nmi & sel_npc_resume}} & npc_r_d1[31:1]));
	rvdffpcie #(.WIDTH(31)) flush_lower_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(tlu_flush_lower_r),
		.din({tlu_flush_path_r[31:1]}),
		.dout({tlu_flush_path_r_d1[31:1]})
	);
	assign dec_tlu_flush_lower_wb = tlu_flush_lower_r_d1;
	assign dec_tlu_flush_lower_r = tlu_flush_lower_r;
	assign dec_tlu_flush_path_r[31:1] = tlu_flush_path_r[31:1];
	assign exc_or_int_valid_r = ((lsu_exc_valid_r | i0_exception_valid_r) | interrupt_valid_r) | (i0_trigger_hit_r & ~trigger_hit_dmode_r);
	rvdffie #(.WIDTH(12)) excinfo_wb_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din({interrupt_valid_r, i0_exception_valid_r, exc_or_int_valid_r, exc_cause_r[4:0], tlu_i0_commit_cmt & ~illegal_r, i0_trigger_hit_r, take_nmi, pause_expired_r}),
		.dout({interrupt_valid_r_d1, i0_exception_valid_r_d1, exc_or_int_valid_r_d1, exc_cause_wb[4:0], i0_valid_wb, trigger_hit_r_d1, take_nmi_r_d1, pause_expired_wb})
	);
	localparam MISA = 12'h301;
	localparam MVENDORID = 12'hf11;
	localparam MARCHID = 12'hf12;
	localparam MIMPID = 12'hf13;
	localparam MHARTID = 12'hf14;
	localparam MSTATUS = 12'h300;
	assign dec_csr_wen_r_mod = (dec_csr_wen_r & ~i0_trigger_hit_r) & ~rfpc_i0_r;
	assign wr_mstatus_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MSTATUS);
	assign set_mie_pmu_fw_halt = ~mpmc_b_ns[1] & fw_halt_req;
	assign mstatus_ns[1:0] = ((((({2 {~wr_mstatus_r & exc_or_int_valid_r}} & {mstatus[MSTATUS_MIE], 1'b0}) | ({2 {wr_mstatus_r & exc_or_int_valid_r}} & {dec_csr_wrdata_r[3], 1'b0})) | ({2 {mret_r & ~exc_or_int_valid_r}} & {1'b1, mstatus[1]})) | ({2 {set_mie_pmu_fw_halt}} & {mstatus[1], 1'b1})) | ({2 {wr_mstatus_r & ~exc_or_int_valid_r}} & {dec_csr_wrdata_r[7], dec_csr_wrdata_r[3]})) | ({2 {((~wr_mstatus_r & ~exc_or_int_valid_r) & ~mret_r) & ~set_mie_pmu_fw_halt}} & mstatus[1:0]);
	assign mstatus_mie_ns = mstatus[MSTATUS_MIE] & (~dcsr_single_step_running_f | dcsr[DCSR_STEPIE]);
	localparam MTVEC = 12'h305;
	assign wr_mtvec_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTVEC);
	assign mtvec_ns[30:0] = {dec_csr_wrdata_r[31:2], dec_csr_wrdata_r[0]};
	rvdffe #(.WIDTH(31)) mtvec_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mtvec_r),
		.din(mtvec_ns[30:0]),
		.dout(mtvec[30:0])
	);
	localparam MIP = 12'h344;
	assign ce_int = (mdccme_ce_req | miccme_ce_req) | mice_ce_req;
	assign mip_ns[5:0] = {ce_int, dec_timer_t0_pulse, dec_timer_t1_pulse, mexintpend, timer_int_sync, soft_int_sync};
	localparam MIE = 12'h304;
	assign wr_mie_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MIE);
	assign mie_ns[5:0] = (wr_mie_r ? {dec_csr_wrdata_r[30:28], dec_csr_wrdata_r[11], dec_csr_wrdata_r[7], dec_csr_wrdata_r[3]} : mie[5:0]);
	rvdff #(.WIDTH(6)) mie_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.din(mie_ns[5:0]),
		.dout(mie[5:0])
	);
	localparam MCYCLEL = 12'hb00;
	assign kill_ebreak_count_r = ebreak_to_debug_mode_r & dcsr[DCSR_STOPC];
	assign wr_mcyclel_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCYCLEL);
	assign mcyclel_cout_in = ~(((kill_ebreak_count_r | (dec_tlu_dbg_halted & dcsr[DCSR_STOPC])) | dec_tlu_pmu_fw_halted) | mcountinhibit[0]);
	assign {mcyclela_cout, mcyclel_inc[7:0]} = mcyclel[7:0] + 8'b00000001;
	assign {mcyclel_cout, mcyclel_inc[31:8]} = mcyclel[31:8] + {23'b00000000000000000000000, mcyclela_cout};
	assign mcyclel_ns[31:0] = (wr_mcyclel_r ? dec_csr_wrdata_r[31:0] : mcyclel_inc[31:0]);
	rvdffe #(.WIDTH(24)) mcyclel_bff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(wr_mcyclel_r | (mcyclela_cout & mcyclel_cout_in)),
		.din(mcyclel_ns[31:8]),
		.dout(mcyclel[31:8])
	);
	rvdffe #(.WIDTH(8)) mcyclel_aff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(wr_mcyclel_r | mcyclel_cout_in),
		.din(mcyclel_ns[7:0]),
		.dout(mcyclel[7:0])
	);
	localparam MCYCLEH = 12'hb80;
	assign wr_mcycleh_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCYCLEH);
	assign mcycleh_inc[31:0] = mcycleh[31:0] + {31'b0000000000000000000000000000000, mcyclel_cout_f};
	assign mcycleh_ns[31:0] = (wr_mcycleh_r ? dec_csr_wrdata_r[31:0] : mcycleh_inc[31:0]);
	rvdffe #(.WIDTH(32)) mcycleh_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(wr_mcycleh_r | mcyclel_cout_f),
		.din(mcycleh_ns[31:0]),
		.dout(mcycleh[31:0])
	);
	localparam MINSTRETL = 12'hb02;
	assign i0_valid_no_ebreak_ecall_r = dec_tlu_i0_valid_r & ~((((ebreak_r | ecall_r) | ebreak_to_debug_mode_r) | illegal_r) | mcountinhibit[2]);
	assign wr_minstretl_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MINSTRETL);
	assign {minstretl_couta, minstretl_inc[7:0]} = minstretl[7:0] + 8'b00000001;
	assign {minstretl_cout, minstretl_inc[31:8]} = minstretl[31:8] + {23'b00000000000000000000000, minstretl_couta};
	assign minstret_enable = (i0_valid_no_ebreak_ecall_r & tlu_i0_commit_cmt) | wr_minstretl_r;
	assign minstretl_cout_ns = ((minstretl_cout & ~wr_minstreth_r) & i0_valid_no_ebreak_ecall_r) & ~dec_tlu_dbg_halted;
	assign minstretl_ns[31:0] = (wr_minstretl_r ? dec_csr_wrdata_r[31:0] : minstretl_inc[31:0]);
	rvdffe #(.WIDTH(24)) minstretl_bff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_minstretl_r | (minstretl_couta & minstret_enable)),
		.din(minstretl_ns[31:8]),
		.dout(minstretl[31:8])
	);
	rvdffe #(.WIDTH(8)) minstretl_aff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(minstret_enable),
		.din(minstretl_ns[7:0]),
		.dout(minstretl[7:0])
	);
	assign minstretl_read[31:0] = minstretl[31:0];
	localparam MINSTRETH = 12'hb82;
	assign wr_minstreth_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MINSTRETH);
	assign minstreth_inc[31:0] = minstreth[31:0] + {31'b0000000000000000000000000000000, minstretl_cout_f};
	assign minstreth_ns[31:0] = (wr_minstreth_r ? dec_csr_wrdata_r[31:0] : minstreth_inc[31:0]);
	rvdffe #(.WIDTH(32)) minstreth_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((minstret_enable_f & minstretl_cout_f) | wr_minstreth_r),
		.din(minstreth_ns[31:0]),
		.dout(minstreth[31:0])
	);
	assign minstreth_read[31:0] = minstreth_inc[31:0];
	localparam MSCRATCH = 12'h340;
	assign wr_mscratch_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MSCRATCH);
	rvdffe #(.WIDTH(32)) mscratch_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mscratch_r),
		.din(dec_csr_wrdata_r[31:0]),
		.dout(mscratch[31:0])
	);
	localparam MEPC = 12'h341;
	assign sel_exu_npc_r = (~dec_tlu_dbg_halted & ~tlu_flush_lower_r_d1) & dec_tlu_i0_valid_r;
	assign sel_flush_npc_r = (~dec_tlu_dbg_halted & tlu_flush_lower_r_d1) & ~dec_tlu_flush_noredir_r_d1;
	assign sel_hold_npc_r = ~sel_exu_npc_r & ~sel_flush_npc_r;
	assign npc_r[31:1] = ((({31 {sel_exu_npc_r}} & exu_npc_r[31:1]) | ({31 {~mpc_reset_run_req & reset_delayed}} & rst_vec[31:1])) | ({31 {sel_flush_npc_r}} & tlu_flush_path_r_d1[31:1])) | ({31 {sel_hold_npc_r}} & npc_r_d1[31:1]);
	rvdffpcie #(.WIDTH(31)) npwbc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((sel_exu_npc_r | sel_flush_npc_r) | reset_delayed),
		.din(npc_r[31:1]),
		.dout(npc_r_d1[31:1])
	);
	assign pc0_valid_r = ~dec_tlu_dbg_halted & dec_tlu_i0_valid_r;
	assign pc_r[31:1] = ({31 {pc0_valid_r}} & dec_tlu_i0_pc_r[31:1]) | ({31 {~pc0_valid_r}} & pc_r_d1[31:1]);
	rvdffpcie #(.WIDTH(31)) pwbc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(pc0_valid_r),
		.din(pc_r[31:1]),
		.dout(pc_r_d1[31:1])
	);
	assign wr_mepc_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEPC);
	assign mepc_ns[31:1] = ((({31 {(i0_exception_valid_r | lsu_exc_valid_r) | mepc_trigger_hit_sel_pc_r}} & pc_r[31:1]) | ({31 {interrupt_valid_r}} & npc_r[31:1])) | ({31 {wr_mepc_r & ~exc_or_int_valid_r}} & dec_csr_wrdata_r[31:1])) | ({31 {~wr_mepc_r & ~exc_or_int_valid_r}} & mepc[31:1]);
	rvdffe #(.WIDTH(31)) mepc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((((i0_exception_valid_r | lsu_exc_valid_r) | mepc_trigger_hit_sel_pc_r) | interrupt_valid_r) | wr_mepc_r),
		.din(mepc_ns[31:1]),
		.dout(mepc[31:1])
	);
	localparam MCAUSE = 12'h342;
	assign wr_mcause_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCAUSE);
	assign mcause_sel_nmi_store = (exc_or_int_valid_r & take_nmi) & nmi_lsu_store_type;
	assign mcause_sel_nmi_load = (exc_or_int_valid_r & take_nmi) & nmi_lsu_load_type;
	assign mcause_sel_nmi_ext = (((exc_or_int_valid_r & take_nmi) & take_ext_int_start_d3) & |lsu_fir_error[1:0]) & ~nmi_int_detected_f;
	assign mcause_fir_error_type[1:0] = {&lsu_fir_error[1:0], lsu_fir_error[1] & ~lsu_fir_error[0]};
	assign mcause_ns[31:0] = ((((({32 {mcause_sel_nmi_store}} & 32'hf0000000) | ({32 {mcause_sel_nmi_load}} & 32'hf0000001)) | ({32 {mcause_sel_nmi_ext}} & {30'b111100000000000000010000000000, mcause_fir_error_type[1:0]})) | ({32 {exc_or_int_valid_r & ~take_nmi}} & {interrupt_valid_r, 26'b00000000000000000000000000, exc_cause_r[4:0]})) | ({32 {wr_mcause_r & ~exc_or_int_valid_r}} & dec_csr_wrdata_r[31:0])) | ({32 {~wr_mcause_r & ~exc_or_int_valid_r}} & mcause[31:0]);
	rvdffe #(.WIDTH(32)) mcause_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(exc_or_int_valid_r | wr_mcause_r),
		.din(mcause_ns[31:0]),
		.dout(mcause[31:0])
	);
	localparam MSCAUSE = 12'h7ff;
	assign wr_mscause_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MSCAUSE);
	assign ifu_mscause[3:0] = (dec_tlu_packet_r[14:13] == 2'b00 ? 4'b1001 : {2'b00, dec_tlu_packet_r[14:13]});
	assign mscause_type[3:0] = ((({4 {lsu_i0_exc_r}} & lsu_error_pkt_r[37:34]) | ({4 {i0_trigger_hit_r}} & 4'b0001)) | ({4 {ebreak_r}} & 4'b0010)) | ({4 {inst_acc_r}} & ifu_mscause[3:0]);
	assign mscause_ns[3:0] = (({4 {exc_or_int_valid_r}} & mscause_type[3:0]) | ({4 {wr_mscause_r & ~exc_or_int_valid_r}} & dec_csr_wrdata_r[3:0])) | ({4 {~wr_mscause_r & ~exc_or_int_valid_r}} & mscause[3:0]);
	rvdff #(.WIDTH(4)) mscause_ff(
		.rst_l(rst_l),
		.clk(e4e5_int_clk),
		.din(mscause_ns[3:0]),
		.dout(mscause[3:0])
	);
	localparam MTVAL = 12'h343;
	assign wr_mtval_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTVAL);
	assign mtval_capture_pc_r = (exc_or_int_valid_r & ((ebreak_r | (inst_acc_r & ~inst_acc_second_r)) | mepc_trigger_hit_sel_pc_r)) & ~take_nmi;
	assign mtval_capture_pc_plus2_r = (exc_or_int_valid_r & (inst_acc_r & inst_acc_second_r)) & ~take_nmi;
	assign mtval_capture_inst_r = (exc_or_int_valid_r & illegal_r) & ~take_nmi;
	assign mtval_capture_lsu_r = (exc_or_int_valid_r & lsu_exc_valid_r) & ~take_nmi;
	assign mtval_clear_r = (((exc_or_int_valid_r & ~mtval_capture_pc_r) & ~mtval_capture_inst_r) & ~mtval_capture_lsu_r) & ~mepc_trigger_hit_sel_pc_r;
	assign mtval_ns[31:0] = ((((({32 {mtval_capture_pc_r}} & {pc_r[31:1], 1'b0}) | ({32 {mtval_capture_pc_plus2_r}} & {pc_r[31:1] + 31'b0000000000000000000000000000001, 1'b0})) | ({32 {mtval_capture_inst_r}} & dec_illegal_inst[31:0])) | ({32 {mtval_capture_lsu_r}} & lsu_error_pkt_addr_r[31:0])) | ({32 {wr_mtval_r & ~interrupt_valid_r}} & dec_csr_wrdata_r[31:0])) | ({32 {((((~take_nmi & ~wr_mtval_r) & ~mtval_capture_pc_r) & ~mtval_capture_inst_r) & ~mtval_clear_r) & ~mtval_capture_lsu_r}} & mtval[31:0]);
	rvdffe #(.WIDTH(32)) mtval_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(tlu_flush_lower_r | wr_mtval_r),
		.din(mtval_ns[31:0]),
		.dout(mtval[31:0])
	);
	localparam MCGC = 12'h7f8;
	assign wr_mcgc_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCGC);
	assign mcgc_ns[9:0] = (wr_mcgc_r ? {~dec_csr_wrdata_r[9], dec_csr_wrdata_r[8:0]} : mcgc_int[9:0]);
	rvdffe #(.WIDTH(10)) mcgc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mcgc_r),
		.din(mcgc_ns[9:0]),
		.dout(mcgc_int[9:0])
	);
	assign mcgc[9:0] = {~mcgc_int[9], mcgc_int[8:0]};
	assign dec_tlu_picio_clk_override = mcgc[9];
	assign dec_tlu_misc_clk_override = mcgc[8];
	assign dec_tlu_dec_clk_override = mcgc[7];
	assign dec_tlu_ifu_clk_override = mcgc[5];
	assign dec_tlu_lsu_clk_override = mcgc[4];
	assign dec_tlu_bus_clk_override = mcgc[3];
	assign dec_tlu_pic_clk_override = mcgc[2];
	assign dec_tlu_dccm_clk_override = mcgc[1];
	assign dec_tlu_icm_clk_override = mcgc[0];
	localparam MFDC = 12'h7f9;
	assign wr_mfdc_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MFDC);
	rvdffe #(.WIDTH(16)) mfdc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mfdc_r),
		.din({mfdc_ns[15:0]}),
		.dout(mfdc_int[15:0])
	);
	generate
		if (pt[2037-:5] == 1) begin : axi4
			assign mfdc_ns[15:0] = {~dec_csr_wrdata_r[18:16], dec_csr_wrdata_r[12], dec_csr_wrdata_r[11:7], ~dec_csr_wrdata_r[6], dec_csr_wrdata_r[5:0]};
			assign mfdc[18:0] = {~mfdc_int[15:13], 3'b000, mfdc_int[12], mfdc_int[11:7], ~mfdc_int[6], mfdc_int[5:0]};
		end
		else begin
			assign mfdc_ns[15:0] = {~dec_csr_wrdata_r[18:16], dec_csr_wrdata_r[12:0]};
			assign mfdc[18:0] = {~mfdc_int[15:13], 3'b000, mfdc_int[12:0]};
		end
	endgenerate
	assign dec_tlu_dma_qos_prty[2:0] = mfdc[18:16];
	assign dec_tlu_trace_disable = mfdc[12];
	assign dec_tlu_external_ldfwd_disable = mfdc[11];
	assign dec_tlu_core_ecc_disable = 1'b1;
	assign dec_tlu_sideeffect_posted_disable = mfdc[6];
	assign dec_tlu_bpred_disable = mfdc[3];
	assign dec_tlu_wb_coalescing_disable = mfdc[2];
	assign dec_tlu_pipelining_disable = mfdc[0];
	assign dec_tlu_wr_pause_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCPC)) & ~interrupt_valid_r) & ~take_ext_int_start;
	localparam MRAC = 12'h7c0;
	assign wr_mrac_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MRAC);
	assign mrac_in[31:0] = {dec_csr_wrdata_r[31], dec_csr_wrdata_r[30] & ~dec_csr_wrdata_r[31], dec_csr_wrdata_r[29], dec_csr_wrdata_r[28] & ~dec_csr_wrdata_r[29], dec_csr_wrdata_r[27], dec_csr_wrdata_r[26] & ~dec_csr_wrdata_r[27], dec_csr_wrdata_r[25], dec_csr_wrdata_r[24] & ~dec_csr_wrdata_r[25], dec_csr_wrdata_r[23], dec_csr_wrdata_r[22] & ~dec_csr_wrdata_r[23], dec_csr_wrdata_r[21], dec_csr_wrdata_r[20] & ~dec_csr_wrdata_r[21], dec_csr_wrdata_r[19], dec_csr_wrdata_r[18] & ~dec_csr_wrdata_r[19], dec_csr_wrdata_r[17], dec_csr_wrdata_r[16] & ~dec_csr_wrdata_r[17], dec_csr_wrdata_r[15], dec_csr_wrdata_r[14] & ~dec_csr_wrdata_r[15], dec_csr_wrdata_r[13], dec_csr_wrdata_r[12] & ~dec_csr_wrdata_r[13], dec_csr_wrdata_r[11], dec_csr_wrdata_r[10] & ~dec_csr_wrdata_r[11], dec_csr_wrdata_r[9], dec_csr_wrdata_r[8] & ~dec_csr_wrdata_r[9], dec_csr_wrdata_r[7], dec_csr_wrdata_r[6] & ~dec_csr_wrdata_r[7], dec_csr_wrdata_r[5], dec_csr_wrdata_r[4] & ~dec_csr_wrdata_r[5], dec_csr_wrdata_r[3], dec_csr_wrdata_r[2] & ~dec_csr_wrdata_r[3], dec_csr_wrdata_r[1], dec_csr_wrdata_r[0] & ~dec_csr_wrdata_r[1]};
	rvdffe #(.WIDTH(32)) mrac_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mrac_r),
		.din(mrac_in[31:0]),
		.dout(mrac[31:0])
	);
	assign dec_tlu_mrac_ff[31:0] = mrac[31:0];
	localparam MDEAU = 12'hbc0;
	assign wr_mdeau_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MDEAU);
	localparam MDSEAC = 12'hfc0;
	assign mdseac_locked_ns = mdseac_en | (mdseac_locked_f & ~wr_mdeau_r);
	assign mdseac_en = ((lsu_imprecise_error_store_any | lsu_imprecise_error_load_any) & ~nmi_int_detected_f) & ~mdseac_locked_f;
	rvdffe #(.WIDTH(32)) mdseac_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(mdseac_en),
		.din(lsu_imprecise_error_addr_any[31:0]),
		.dout(mdseac[31:0])
	);
	localparam MPMC = 12'h7c6;
	assign wr_mpmc_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MPMC);
	assign fw_halt_req = ((wr_mpmc_r & dec_csr_wrdata_r[0]) & ~internal_dbg_halt_mode_f2) & ~ext_int_freeze_d1;
	assign fw_halted_ns = (fw_halt_req | fw_halted) & ~set_mie_pmu_fw_halt;
	assign mpmc_b_ns[1] = (wr_mpmc_r ? ~dec_csr_wrdata_r[1] : ~mpmc[1]);
	rvdff #(.WIDTH(1)) mpmc_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.din(mpmc_b_ns[1]),
		.dout(mpmc_b[1])
	);
	assign mpmc[1] = ~mpmc_b[1];
	localparam MICECT = 12'h7f0;
	assign csr_sat[31:27] = (dec_csr_wrdata_r[31:27] > 5'd26 ? 5'd26 : dec_csr_wrdata_r[31:27]);
	assign wr_micect_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MICECT);
	assign micect_inc[26:0] = micect[26:0] + {26'b00000000000000000000000000, ic_perr_r};
	assign micect_ns = (wr_micect_r ? {csr_sat[31:27], dec_csr_wrdata_r[26:0]} : {micect[31:27], micect_inc[26:0]});
	rvdffe #(.WIDTH(32)) micect_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_micect_r | ic_perr_r),
		.din(micect_ns[31:0]),
		.dout(micect[31:0])
	);
	assign mice_ce_req = |({32'hffffffff << micect[31:27]} & {5'b00000, micect[26:0]});
	localparam MICCMECT = 12'h7f1;
	assign wr_miccmect_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MICCMECT);
	assign miccmect_inc[26:0] = miccmect[26:0] + {26'b00000000000000000000000000, iccm_sbecc_r | iccm_dma_sb_error};
	assign miccmect_ns = (wr_miccmect_r ? {csr_sat[31:27], dec_csr_wrdata_r[26:0]} : {miccmect[31:27], miccmect_inc[26:0]});
	rvdffe #(.WIDTH(32)) miccmect_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en((wr_miccmect_r | iccm_sbecc_r) | iccm_dma_sb_error),
		.din(miccmect_ns[31:0]),
		.dout(miccmect[31:0])
	);
	assign miccme_ce_req = |({32'hffffffff << miccmect[31:27]} & {5'b00000, miccmect[26:0]});
	localparam MDCCMECT = 12'h7f2;
	assign wr_mdccmect_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MDCCMECT);
	assign mdccmect_inc[26:0] = mdccmect[26:0] + {26'b00000000000000000000000000, lsu_single_ecc_error_r_d1};
	assign mdccmect_ns = (wr_mdccmect_r ? {csr_sat[31:27], dec_csr_wrdata_r[26:0]} : {mdccmect[31:27], mdccmect_inc[26:0]});
	rvdffe #(.WIDTH(32)) mdccmect_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(wr_mdccmect_r | lsu_single_ecc_error_r_d1),
		.din(mdccmect_ns[31:0]),
		.dout(mdccmect[31:0])
	);
	assign mdccme_ce_req = |({32'hffffffff << mdccmect[31:27]} & {5'b00000, mdccmect[26:0]});
	localparam MFDHT = 12'h7ce;
	assign wr_mfdht_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MFDHT);
	assign mfdht_ns[5:0] = (wr_mfdht_r ? dec_csr_wrdata_r[5:0] : mfdht[5:0]);
	rvdffs #(.WIDTH(6)) mfdht_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.en(wr_mfdht_r),
		.din(mfdht_ns[5:0]),
		.dout(mfdht[5:0])
	);
	localparam MFDHS = 12'h7cf;
	assign wr_mfdhs_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MFDHS);
	assign mfdhs_ns[1:0] = (wr_mfdhs_r ? dec_csr_wrdata_r[1:0] : (dbg_tlu_halted & ~dbg_tlu_halted_f ? {~lsu_idle_any_f, ~ifu_miss_state_idle_f} : mfdhs[1:0]));
	rvdffs #(.WIDTH(2)) mfdhs_ff(
		.rst_l(rst_l),
		.clk(free_clk),
		.en(wr_mfdhs_r | dbg_tlu_halted),
		.din(mfdhs_ns[1:0]),
		.dout(mfdhs[1:0])
	);
	assign force_halt_ctr[31:0] = (debug_halt_req_f ? force_halt_ctr_f[31:0] + 32'b00000000000000000000000000000001 : (dbg_tlu_halted_f ? 32'b00000000000000000000000000000000 : force_halt_ctr_f[31:0]));
	rvdffe #(.WIDTH(32)) forcehaltctr_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(mfdht[0]),
		.din(force_halt_ctr[31:0]),
		.dout(force_halt_ctr_f[31:0])
	);
	assign force_halt = mfdht[0] & |(force_halt_ctr_f[31:0] & (32'hffffffff << mfdht[5:1]));
	localparam MEIVT = 12'hbc8;
	assign wr_meivt_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEIVT);
	rvdffe #(.WIDTH(22)) meivt_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_meivt_r),
		.din(dec_csr_wrdata_r[31:10]),
		.dout(meivt[31:10])
	);
	localparam MEIHAP = 12'hfc8;
	assign wr_meihap_r = wr_meicpct_r;
	rvdffe #(.WIDTH(8)) meihap_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_meihap_r),
		.din(pic_claimid[7:0]),
		.dout(meihap[9:2])
	);
	assign dec_tlu_meihap[31:2] = {meivt[31:10], meihap[9:2]};
	localparam MEICURPL = 12'hbcc;
	assign wr_meicurpl_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEICURPL);
	assign meicurpl_ns[3:0] = (wr_meicurpl_r ? dec_csr_wrdata_r[3:0] : meicurpl[3:0]);
	rvdff #(.WIDTH(4)) meicurpl_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.din(meicurpl_ns[3:0]),
		.dout(meicurpl[3:0])
	);
	assign dec_tlu_meicurpl[3:0] = meicurpl[3:0];
	localparam MEICIDPL = 12'hbcb;
	assign wr_meicidpl_r = (dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEICIDPL)) | take_ext_int_start;
	assign meicidpl_ns[3:0] = (wr_meicpct_r ? pic_pl[3:0] : (wr_meicidpl_r ? dec_csr_wrdata_r[3:0] : meicidpl[3:0]));
	localparam MEICPCT = 12'hbca;
	assign wr_meicpct_r = (dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEICPCT)) | take_ext_int_start;
	localparam MEIPT = 12'hbc9;
	assign wr_meipt_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MEIPT);
	assign meipt_ns[3:0] = (wr_meipt_r ? dec_csr_wrdata_r[3:0] : meipt[3:0]);
	rvdff #(.WIDTH(4)) meipt_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.din(meipt_ns[3:0]),
		.dout(meipt[3:0])
	);
	assign dec_tlu_meipt[3:0] = meipt[3:0];
	localparam DCSR = 12'h7b0;
	assign trigger_hit_for_dscr_cause_r_d1 = trigger_hit_dmode_r_d1 | (trigger_hit_r_d1 & dcsr_single_step_done_f);
	assign dcsr_cause[8:6] = ((({3 {((dcsr_single_step_done_f & ~ebreak_to_debug_mode_r_d1) & ~trigger_hit_for_dscr_cause_r_d1) & ~debug_halt_req}} & 3'b100) | ({3 {(debug_halt_req & ~ebreak_to_debug_mode_r_d1) & ~trigger_hit_for_dscr_cause_r_d1}} & 3'b011)) | ({3 {ebreak_to_debug_mode_r_d1 & ~trigger_hit_for_dscr_cause_r_d1}} & 3'b001)) | ({3 {trigger_hit_for_dscr_cause_r_d1}} & 3'b010);
	assign wr_dcsr_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DCSR);
	assign dcsr_cause_upgradeable = internal_dbg_halt_mode_f & (dcsr[8:6] == 3'b011);
	assign enter_debug_halt_req_le = enter_debug_halt_req & (~dbg_tlu_halted | dcsr_cause_upgradeable);
	assign nmi_in_debug_mode = nmi_int_detected_f & internal_dbg_halt_mode_f;
	assign dcsr_ns[15:2] = (enter_debug_halt_req_le ? {dcsr[15:9], dcsr_cause[8:6], dcsr[5:2]} : (wr_dcsr_r ? {dec_csr_wrdata_r[15], 3'b000, dec_csr_wrdata_r[11:10], 1'b0, dcsr[8:6], 2'b00, nmi_in_debug_mode | dcsr[3], dec_csr_wrdata_r[2]} : {dcsr[15:4], nmi_in_debug_mode, dcsr[2]}));
	rvdffe #(.WIDTH(14)) dcsr_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(((enter_debug_halt_req_le | wr_dcsr_r) | internal_dbg_halt_mode) | take_nmi),
		.din(dcsr_ns[15:2]),
		.dout(dcsr[15:2])
	);
	localparam DPC = 12'h7b1;
	assign wr_dpc_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DPC);
	assign dpc_capture_npc = (dbg_tlu_halted & ~dbg_tlu_halted_f) & ~request_debug_mode_done;
	assign dpc_capture_pc = request_debug_mode_r;
	assign dpc_ns[31:1] = (({31 {(~dpc_capture_pc & ~dpc_capture_npc) & wr_dpc_r}} & dec_csr_wrdata_r[31:1]) | ({31 {dpc_capture_pc}} & pc_r[31:1])) | ({31 {~dpc_capture_pc & dpc_capture_npc}} & npc_r[31:1]);
	rvdffe #(.WIDTH(31)) dpc_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((wr_dpc_r | dpc_capture_pc) | dpc_capture_npc),
		.din(dpc_ns[31:1]),
		.dout(dpc[31:1])
	);
	localparam DICAWICS = 12'h7c8;
	assign dicawics_ns[16:0] = {dec_csr_wrdata_r[24], dec_csr_wrdata_r[21:20], dec_csr_wrdata_r[16:3]};
	assign wr_dicawics_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAWICS);
	rvdffe #(.WIDTH(17)) dicawics_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_dicawics_r),
		.din(dicawics_ns[16:0]),
		.dout(dicawics[16:0])
	);
	localparam DICAD0 = 12'h7c9;
	assign dicad0_ns[31:0] = (wr_dicad0_r ? dec_csr_wrdata_r[31:0] : ifu_ic_debug_rd_data[31:0]);
	assign wr_dicad0_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAD0);
	rvdffe #(.WIDTH(32)) dicad0_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_dicad0_r | ifu_ic_debug_rd_data_valid),
		.din(dicad0_ns[31:0]),
		.dout(dicad0[31:0])
	);
	localparam DICAD0H = 12'h7cc;
	assign dicad0h_ns[31:0] = (wr_dicad0h_r ? dec_csr_wrdata_r[31:0] : ifu_ic_debug_rd_data[63:32]);
	assign wr_dicad0h_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAD0H);
	rvdffe #(.WIDTH(32)) dicad0h_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_dicad0h_r | ifu_ic_debug_rd_data_valid),
		.din(dicad0h_ns[31:0]),
		.dout(dicad0h[31:0])
	);
	generate
		if (pt[1125-:5] == 1) begin
			localparam DICAD1 = 12'h7ca;
			assign dicad1_ns[6:0] = (wr_dicad1_r ? dec_csr_wrdata_r[6:0] : ifu_ic_debug_rd_data[70:64]);
			assign wr_dicad1_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAD1);
			rvdffe #(
				.WIDTH(7),
				.OVERRIDE(1)
			) dicad1_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(wr_dicad1_r | ifu_ic_debug_rd_data_valid),
				.din(dicad1_ns[6:0]),
				.dout(dicad1_raw[6:0])
			);
			assign dicad1[31:0] = {25'b0000000000000000000000000, dicad1_raw[6:0]};
		end
		else begin
			localparam DICAD1 = 12'h7ca;
			assign dicad1_ns[3:0] = (wr_dicad1_r ? dec_csr_wrdata_r[3:0] : ifu_ic_debug_rd_data[67:64]);
			assign wr_dicad1_r = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAD1);
			rvdffs #(.WIDTH(4)) dicad1_ff(
				.rst_l(rst_l),
				.clk(free_clk),
				.en(wr_dicad1_r | ifu_ic_debug_rd_data_valid),
				.din(dicad1_ns[3:0]),
				.dout(dicad1_raw[3:0])
			);
			assign dicad1[31:0] = {28'b0000000000000000000000000000, dicad1_raw[3:0]};
		end
	endgenerate
	localparam DICAGO = 12'h7cb;
	generate
		if (pt[1125-:5] == 1) begin
			assign dec_tlu_ic_diag_pkt[89:19] = {dicad1[6:0], dicad0h[31:0], dicad0[31:0]};
		end
		else assign dec_tlu_ic_diag_pkt[89:19] = {3'b000, dicad1[3:0], dicad0h[31:0], dicad0[31:0]};
	endgenerate
	assign dec_tlu_ic_diag_pkt[18:2] = dicawics[16:0];
	assign icache_rd_valid = (((allow_dbg_halt_csr_write & dec_csr_any_unq_d) & dec_i0_decode_d) & ~dec_csr_wen_unq_d) & (dec_csr_rdaddr_d[11:0] == DICAGO);
	assign icache_wr_valid = (allow_dbg_halt_csr_write & dec_csr_wen_r_mod) & (dec_csr_wraddr_r[11:0] == DICAGO);
	assign dec_tlu_ic_diag_pkt[1] = icache_rd_valid_f;
	assign dec_tlu_ic_diag_pkt[0] = icache_wr_valid_f;
	localparam MTSEL = 12'h7a0;
	assign wr_mtsel_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTSEL);
	assign mtsel_ns[1:0] = (wr_mtsel_r ? {dec_csr_wrdata_r[1:0]} : mtsel[1:0]);
	rvdff #(.WIDTH(2)) mtsel_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.din(mtsel_ns[1:0]),
		.dout(mtsel[1:0])
	);
	localparam MTDATA1 = 12'h7a1;
	assign tdata_load = dec_csr_wrdata_r[0] & ~dec_csr_wrdata_r[19];
	assign tdata_opcode = dec_csr_wrdata_r[2] & ~dec_csr_wrdata_r[19];
	assign tdata_action = (dec_csr_wrdata_r[27] & dbg_tlu_halted_f) & dec_csr_wrdata_r[12];
	assign tdata_chain = (mtsel[0] ? 1'b0 : (mtsel[1] ? dec_csr_wrdata_r[11] & ~(mtdata1_t3[MTDATA1_DMODE] & ~dec_csr_wrdata_r[27]) : dec_csr_wrdata_r[11] & ~(mtdata1_t1[MTDATA1_DMODE] & ~dec_csr_wrdata_r[27])));
	assign tdata_kill_write = (mtsel[1] ? dec_csr_wrdata_r[27] & (~mtdata1_t2[MTDATA1_DMODE] & mtdata1_t2[MTDATA1_CHAIN]) : dec_csr_wrdata_r[27] & (~mtdata1_t0[MTDATA1_DMODE] & mtdata1_t0[MTDATA1_CHAIN]));
	assign tdata_wrdata_r[9:0] = {dec_csr_wrdata_r[27] & dbg_tlu_halted_f, dec_csr_wrdata_r[20:19], tdata_action, tdata_chain, dec_csr_wrdata_r[7:6], tdata_opcode, dec_csr_wrdata_r[1], tdata_load};
	assign wr_mtdata1_t0_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA1)) & (mtsel[1:0] == 2'b00)) & (~mtdata1_t0[MTDATA1_DMODE] | dbg_tlu_halted_f);
	assign mtdata1_t0_ns[9:0] = (wr_mtdata1_t0_r ? tdata_wrdata_r[9:0] : {mtdata1_t0[9], update_hit_bit_r[0] | mtdata1_t0[8], mtdata1_t0[7:0]});
	assign wr_mtdata1_t1_r = (((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA1)) & (mtsel[1:0] == 2'b01)) & (~mtdata1_t1[MTDATA1_DMODE] | dbg_tlu_halted_f)) & ~tdata_kill_write;
	assign mtdata1_t1_ns[9:0] = (wr_mtdata1_t1_r ? tdata_wrdata_r[9:0] : {mtdata1_t1[9], update_hit_bit_r[1] | mtdata1_t1[8], mtdata1_t1[7:0]});
	assign wr_mtdata1_t2_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA1)) & (mtsel[1:0] == 2'b10)) & (~mtdata1_t2[MTDATA1_DMODE] | dbg_tlu_halted_f);
	assign mtdata1_t2_ns[9:0] = (wr_mtdata1_t2_r ? tdata_wrdata_r[9:0] : {mtdata1_t2[9], update_hit_bit_r[2] | mtdata1_t2[8], mtdata1_t2[7:0]});
	assign wr_mtdata1_t3_r = (((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA1)) & (mtsel[1:0] == 2'b11)) & (~mtdata1_t3[MTDATA1_DMODE] | dbg_tlu_halted_f)) & ~tdata_kill_write;
	assign mtdata1_t3_ns[9:0] = (wr_mtdata1_t3_r ? tdata_wrdata_r[9:0] : {mtdata1_t3[9], update_hit_bit_r[3] | mtdata1_t3[8], mtdata1_t3[7:0]});
	rvdffe #(.WIDTH(10)) mtdata1_t0_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(trigger_enabled[0] | wr_mtdata1_t0_r),
		.din(mtdata1_t0_ns[9:0]),
		.dout(mtdata1_t0[9:0])
	);
	rvdffe #(.WIDTH(10)) mtdata1_t1_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(trigger_enabled[1] | wr_mtdata1_t1_r),
		.din(mtdata1_t1_ns[9:0]),
		.dout(mtdata1_t1[9:0])
	);
	rvdffe #(.WIDTH(10)) mtdata1_t2_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(trigger_enabled[2] | wr_mtdata1_t2_r),
		.din(mtdata1_t2_ns[9:0]),
		.dout(mtdata1_t2[9:0])
	);
	rvdffe #(.WIDTH(10)) mtdata1_t3_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(trigger_enabled[3] | wr_mtdata1_t3_r),
		.din(mtdata1_t3_ns[9:0]),
		.dout(mtdata1_t3[9:0])
	);
	assign mtdata1_tsel_out[31:0] = ((({32 {mtsel[1:0] == 2'b00}} & {4'h2, mtdata1_t0[9], 6'b011111, mtdata1_t0[8:7], 6'b000000, mtdata1_t0[6:5], 3'b000, mtdata1_t0[4:3], 3'b000, mtdata1_t0[2:0]}) | ({32 {mtsel[1:0] == 2'b01}} & {4'h2, mtdata1_t1[9], 6'b011111, mtdata1_t1[8:7], 6'b000000, mtdata1_t1[6:5], 3'b000, mtdata1_t1[4:3], 3'b000, mtdata1_t1[2:0]})) | ({32 {mtsel[1:0] == 2'b10}} & {4'h2, mtdata1_t2[9], 6'b011111, mtdata1_t2[8:7], 6'b000000, mtdata1_t2[6:5], 3'b000, mtdata1_t2[4:3], 3'b000, mtdata1_t2[2:0]})) | ({32 {mtsel[1:0] == 2'b11}} & {4'h2, mtdata1_t3[9], 6'b011111, mtdata1_t3[8:7], 6'b000000, mtdata1_t3[6:5], 3'b000, mtdata1_t3[4:3], 3'b000, mtdata1_t3[2:0]});
	assign trigger_pkt_any[37] = mtdata1_t0[MTDATA1_SEL];
	assign trigger_pkt_any[36] = mtdata1_t0[MTDATA1_MATCH];
	assign trigger_pkt_any[35] = mtdata1_t0[MTDATA1_ST];
	assign trigger_pkt_any[34] = mtdata1_t0[MTDATA1_LD];
	assign trigger_pkt_any[33] = mtdata1_t0[MTDATA1_EXE];
	assign trigger_pkt_any[32] = mtdata1_t0[MTDATA1_M_ENABLED];
	assign trigger_pkt_any[75] = mtdata1_t1[MTDATA1_SEL];
	assign trigger_pkt_any[74] = mtdata1_t1[MTDATA1_MATCH];
	assign trigger_pkt_any[73] = mtdata1_t1[MTDATA1_ST];
	assign trigger_pkt_any[72] = mtdata1_t1[MTDATA1_LD];
	assign trigger_pkt_any[71] = mtdata1_t1[MTDATA1_EXE];
	assign trigger_pkt_any[70] = mtdata1_t1[MTDATA1_M_ENABLED];
	assign trigger_pkt_any[113] = mtdata1_t2[MTDATA1_SEL];
	assign trigger_pkt_any[112] = mtdata1_t2[MTDATA1_MATCH];
	assign trigger_pkt_any[111] = mtdata1_t2[MTDATA1_ST];
	assign trigger_pkt_any[110] = mtdata1_t2[MTDATA1_LD];
	assign trigger_pkt_any[109] = mtdata1_t2[MTDATA1_EXE];
	assign trigger_pkt_any[108] = mtdata1_t2[MTDATA1_M_ENABLED];
	assign trigger_pkt_any[151] = mtdata1_t3[MTDATA1_SEL];
	assign trigger_pkt_any[150] = mtdata1_t3[MTDATA1_MATCH];
	assign trigger_pkt_any[149] = mtdata1_t3[MTDATA1_ST];
	assign trigger_pkt_any[148] = mtdata1_t3[MTDATA1_LD];
	assign trigger_pkt_any[147] = mtdata1_t3[MTDATA1_EXE];
	assign trigger_pkt_any[146] = mtdata1_t3[MTDATA1_M_ENABLED];
	localparam MTDATA2 = 12'h7a2;
	assign wr_mtdata2_t0_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA2)) & (mtsel[1:0] == 2'b00)) & (~mtdata1_t0[MTDATA1_DMODE] | dbg_tlu_halted_f);
	assign wr_mtdata2_t1_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA2)) & (mtsel[1:0] == 2'b01)) & (~mtdata1_t1[MTDATA1_DMODE] | dbg_tlu_halted_f);
	assign wr_mtdata2_t2_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA2)) & (mtsel[1:0] == 2'b10)) & (~mtdata1_t2[MTDATA1_DMODE] | dbg_tlu_halted_f);
	assign wr_mtdata2_t3_r = ((dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MTDATA2)) & (mtsel[1:0] == 2'b11)) & (~mtdata1_t3[MTDATA1_DMODE] | dbg_tlu_halted_f);
	rvdffe #(.WIDTH(32)) mtdata2_t0_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mtdata2_t0_r),
		.din(dec_csr_wrdata_r[31:0]),
		.dout(mtdata2_t0[31:0])
	);
	rvdffe #(.WIDTH(32)) mtdata2_t1_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mtdata2_t1_r),
		.din(dec_csr_wrdata_r[31:0]),
		.dout(mtdata2_t1[31:0])
	);
	rvdffe #(.WIDTH(32)) mtdata2_t2_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mtdata2_t2_r),
		.din(dec_csr_wrdata_r[31:0]),
		.dout(mtdata2_t2[31:0])
	);
	rvdffe #(.WIDTH(32)) mtdata2_t3_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mtdata2_t3_r),
		.din(dec_csr_wrdata_r[31:0]),
		.dout(mtdata2_t3[31:0])
	);
	assign mtdata2_tsel_out[31:0] = ((({32 {mtsel[1:0] == 2'b00}} & mtdata2_t0[31:0]) | ({32 {mtsel[1:0] == 2'b01}} & mtdata2_t1[31:0])) | ({32 {mtsel[1:0] == 2'b10}} & mtdata2_t2[31:0])) | ({32 {mtsel[1:0] == 2'b11}} & mtdata2_t3[31:0]);
	assign trigger_pkt_any[31-:32] = mtdata2_t0[31:0];
	assign trigger_pkt_any[69-:32] = mtdata2_t1[31:0];
	assign trigger_pkt_any[107-:32] = mtdata2_t2[31:0];
	assign trigger_pkt_any[145-:32] = mtdata2_t3[31:0];
	localparam MHPME_NOEVENT = 10'd0;
	localparam MHPME_CLK_ACTIVE = 10'd1;
	localparam MHPME_ICACHE_HIT = 10'd2;
	localparam MHPME_ICACHE_MISS = 10'd3;
	localparam MHPME_INST_COMMIT = 10'd4;
	localparam MHPME_INST_COMMIT_16B = 10'd5;
	localparam MHPME_INST_COMMIT_32B = 10'd6;
	localparam MHPME_INST_ALIGNED = 10'd7;
	localparam MHPME_INST_DECODED = 10'd8;
	localparam MHPME_INST_MUL = 10'd9;
	localparam MHPME_INST_DIV = 10'd10;
	localparam MHPME_INST_LOAD = 10'd11;
	localparam MHPME_INST_STORE = 10'd12;
	localparam MHPME_INST_MALOAD = 10'd13;
	localparam MHPME_INST_MASTORE = 10'd14;
	localparam MHPME_INST_ALU = 10'd15;
	localparam MHPME_INST_CSRREAD = 10'd16;
	localparam MHPME_INST_CSRRW = 10'd17;
	localparam MHPME_INST_CSRWRITE = 10'd18;
	localparam MHPME_INST_EBREAK = 10'd19;
	localparam MHPME_INST_ECALL = 10'd20;
	localparam MHPME_INST_FENCE = 10'd21;
	localparam MHPME_INST_FENCEI = 10'd22;
	localparam MHPME_INST_MRET = 10'd23;
	localparam MHPME_INST_BRANCH = 10'd24;
	localparam MHPME_BRANCH_MP = 10'd25;
	localparam MHPME_BRANCH_TAKEN = 10'd26;
	localparam MHPME_BRANCH_NOTP = 10'd27;
	localparam MHPME_FETCH_STALL = 10'd28;
	localparam MHPME_DECODE_STALL = 10'd30;
	localparam MHPME_POSTSYNC_STALL = 10'd31;
	localparam MHPME_PRESYNC_STALL = 10'd32;
	localparam MHPME_LSU_SB_WB_STALL = 10'd34;
	localparam MHPME_DMA_DCCM_STALL = 10'd35;
	localparam MHPME_DMA_ICCM_STALL = 10'd36;
	localparam MHPME_EXC_TAKEN = 10'd37;
	localparam MHPME_TIMER_INT_TAKEN = 10'd38;
	localparam MHPME_EXT_INT_TAKEN = 10'd39;
	localparam MHPME_FLUSH_LOWER = 10'd40;
	localparam MHPME_BR_ERROR = 10'd41;
	localparam MHPME_IBUS_TRANS = 10'd42;
	localparam MHPME_DBUS_TRANS = 10'd43;
	localparam MHPME_DBUS_MA_TRANS = 10'd44;
	localparam MHPME_IBUS_ERROR = 10'd45;
	localparam MHPME_DBUS_ERROR = 10'd46;
	localparam MHPME_IBUS_STALL = 10'd47;
	localparam MHPME_DBUS_STALL = 10'd48;
	localparam MHPME_INT_DISABLED = 10'd49;
	localparam MHPME_INT_STALLED = 10'd50;
	localparam MHPME_INST_BITMANIP = 10'd54;
	localparam MHPME_DBUS_LOAD = 10'd55;
	localparam MHPME_DBUS_STORE = 10'd56;
	localparam MHPME_SLEEP_CYC = 10'd512;
	localparam MHPME_DMA_READ_ALL = 10'd513;
	localparam MHPME_DMA_WRITE_ALL = 10'd514;
	localparam MHPME_DMA_READ_DCCM = 10'd515;
	localparam MHPME_DMA_WRITE_DCCM = 10'd516;
	assign mhpme_vec[9-:10] = mhpme3[9:0];
	assign mhpme_vec[19-:10] = mhpme4[9:0];
	assign mhpme_vec[29-:10] = mhpme5[9:0];
	assign mhpme_vec[39-:10] = mhpme6[9:0];
	assign pmu_i0_itype_qual[3:0] = dec_tlu_packet_r[3:0] & {4 {tlu_i0_commit_cmt}};
	localparam [3:0] eb1_pkg_ALU = 4'b0100;
	localparam [3:0] eb1_pkg_BITMANIPU = 4'b1111;
	localparam [3:0] eb1_pkg_CONDBR = 4'b1101;
	localparam [3:0] eb1_pkg_CSRREAD = 4'b0101;
	localparam [3:0] eb1_pkg_CSRRW = 4'b0111;
	localparam [3:0] eb1_pkg_CSRWRITE = 4'b0110;
	localparam [3:0] eb1_pkg_FENCE = 4'b1010;
	localparam [3:0] eb1_pkg_FENCEI = 4'b1011;
	localparam [3:0] eb1_pkg_JAL = 4'b1110;
	localparam [3:0] eb1_pkg_LOAD = 4'b0010;
	localparam [3:0] eb1_pkg_MUL = 4'b0001;
	localparam [3:0] eb1_pkg_STORE = 4'b0011;
	generate
		genvar i;
		for (i = 0; i < 4; i = i + 1) assign mhpmc_inc_r[i] = {~mcountinhibit[i + 3]} & ((((((((((((((((((((((((((((((((((((((((((((((((((((((((({mhpme_vec[(i * 10) + 9-:10] == MHPME_CLK_ACTIVE} & 1'b1) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_ICACHE_HIT} & {ifu_pmu_ic_hit})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_ICACHE_MISS} & {ifu_pmu_ic_miss})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_COMMIT} & {tlu_i0_commit_cmt & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_COMMIT_16B} & {(tlu_i0_commit_cmt & ~exu_pmu_i0_pc4) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_COMMIT_32B} & {(tlu_i0_commit_cmt & exu_pmu_i0_pc4) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_ALIGNED} & ifu_pmu_instr_aligned)) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_DECODED} & dec_pmu_instr_decoded)) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DECODE_STALL} & {dec_pmu_decode_stall})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_MUL} & {pmu_i0_itype_qual == eb1_pkg_MUL})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_DIV} & {(dec_tlu_packet_r[6] & tlu_i0_commit_cmt) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_LOAD} & {pmu_i0_itype_qual == eb1_pkg_LOAD})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_STORE} & {pmu_i0_itype_qual == eb1_pkg_STORE})) | (({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_MALOAD} & {pmu_i0_itype_qual == eb1_pkg_LOAD}) & {dec_tlu_packet_r[4]})) | (({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_MASTORE} & {pmu_i0_itype_qual == eb1_pkg_STORE}) & {dec_tlu_packet_r[4]})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_ALU} & {pmu_i0_itype_qual == eb1_pkg_ALU})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_CSRREAD} & {pmu_i0_itype_qual == eb1_pkg_CSRREAD})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_CSRWRITE} & {pmu_i0_itype_qual == eb1_pkg_CSRWRITE})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_CSRRW} & {pmu_i0_itype_qual == eb1_pkg_CSRRW})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_EBREAK} & {pmu_i0_itype_qual == eb1_pkg_EBREAK})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_ECALL} & {pmu_i0_itype_qual == eb1_pkg_ECALL})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_FENCE} & {pmu_i0_itype_qual == eb1_pkg_FENCE})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_FENCEI} & {pmu_i0_itype_qual == eb1_pkg_FENCEI})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_MRET} & {pmu_i0_itype_qual == eb1_pkg_MRET})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_BRANCH} & {(pmu_i0_itype_qual == eb1_pkg_CONDBR) | (pmu_i0_itype_qual == eb1_pkg_JAL)})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_BRANCH_MP} & {(exu_pmu_i0_br_misp & tlu_i0_commit_cmt) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_BRANCH_TAKEN} & {(exu_pmu_i0_br_ataken & tlu_i0_commit_cmt) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_BRANCH_NOTP} & {(dec_tlu_packet_r[7] & tlu_i0_commit_cmt) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_FETCH_STALL} & {ifu_pmu_fetch_stall})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DECODE_STALL} & {dec_pmu_decode_stall})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_POSTSYNC_STALL} & {dec_pmu_postsync_stall})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_PRESYNC_STALL} & {dec_pmu_presync_stall})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_LSU_SB_WB_STALL} & {lsu_store_stall_any})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_DCCM_STALL} & {dma_dccm_stall_any})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_ICCM_STALL} & {dma_iccm_stall_any})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_EXC_TAKEN} & {(i0_exception_valid_r | i0_trigger_hit_r) | lsu_exc_valid_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_TIMER_INT_TAKEN} & {(take_timer_int | take_int_timer0_int) | take_int_timer1_int})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_EXT_INT_TAKEN} & {take_ext_int})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_FLUSH_LOWER} & {tlu_flush_lower_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_BR_ERROR} & {(dec_tlu_br0_error_r | dec_tlu_br0_start_error_r) & rfpc_i0_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_IBUS_TRANS} & {ifu_pmu_bus_trxn})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_TRANS} & {lsu_pmu_bus_trxn})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_MA_TRANS} & {lsu_pmu_bus_misaligned})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_IBUS_ERROR} & {ifu_pmu_bus_error})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_ERROR} & {lsu_pmu_bus_error})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_IBUS_STALL} & {ifu_pmu_bus_busy})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_STALL} & {lsu_pmu_bus_busy})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INT_DISABLED} & {~mstatus[MSTATUS_MIE]})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INT_STALLED} & {~mstatus[MSTATUS_MIE] & |(mip[5:0] & mie[5:0])})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_INST_BITMANIP} & {pmu_i0_itype_qual == eb1_pkg_BITMANIPU})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_LOAD} & {(tlu_i0_commit_cmt & lsu_pmu_load_external_r) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DBUS_STORE} & {(tlu_i0_commit_cmt & lsu_pmu_store_external_r) & ~illegal_r})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_SLEEP_CYC} & {dec_tlu_pmu_fw_halted})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_READ_ALL} & {dma_pmu_any_read})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_WRITE_ALL} & {dma_pmu_any_write})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_READ_DCCM} & {dma_pmu_dccm_read})) | ({mhpme_vec[(i * 10) + 9-:10] == MHPME_DMA_WRITE_DCCM} & {dma_pmu_dccm_write}));
	endgenerate
	generate
		if (pt[1227-:5]) begin
			rvdffie #(.WIDTH(31)) mstatus_ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(free_l2clk),
				.din({mdseac_locked_ns, lsu_single_ecc_error_r, lsu_exc_valid_r, lsu_i0_exc_r, take_ext_int_start, take_ext_int_start_d1, take_ext_int_start_d2, ext_int_freeze, mip_ns[5:0], (mcyclel_cout & ~wr_mcycleh_r) & mcyclel_cout_in, minstret_enable, minstretl_cout_ns, fw_halted_ns, meicidpl_ns[3:0], icache_rd_valid, icache_wr_valid, mhpmc_inc_r[3:0], perfcnt_halted, mstatus_ns[1:0]}),
				.dout({mdseac_locked_f, lsu_single_ecc_error_r_d1, lsu_exc_valid_r_d1, lsu_i0_exc_r_d1, take_ext_int_start_d1, take_ext_int_start_d2, take_ext_int_start_d3, ext_int_freeze_d1, mip[5:0], mcyclel_cout_f, minstret_enable_f, minstretl_cout_f, fw_halted, meicidpl[3:0], icache_rd_valid_f, icache_wr_valid_f, mhpmc_inc_r_d1[3:0], perfcnt_halted_d1, mstatus[1:0]})
			);
		end
		else rvdffie #(.WIDTH(27)) mstatus_ff(
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.clk(free_l2clk),
			.din({mdseac_locked_ns, lsu_single_ecc_error_r, lsu_exc_valid_r, lsu_i0_exc_r, mip_ns[5:0], (mcyclel_cout & ~wr_mcycleh_r) & mcyclel_cout_in, minstret_enable, minstretl_cout_ns, fw_halted_ns, meicidpl_ns[3:0], icache_rd_valid, icache_wr_valid, mhpmc_inc_r[3:0], perfcnt_halted, mstatus_ns[1:0]}),
			.dout({mdseac_locked_f, lsu_single_ecc_error_r_d1, lsu_exc_valid_r_d1, lsu_i0_exc_r_d1, mip[5:0], mcyclel_cout_f, minstret_enable_f, minstretl_cout_f, fw_halted, meicidpl[3:0], icache_rd_valid_f, icache_wr_valid_f, mhpmc_inc_r_d1[3:0], perfcnt_halted_d1, mstatus[1:0]})
		);
	endgenerate
	assign perfcnt_halted = (dec_tlu_dbg_halted & dcsr[DCSR_STOPC]) | dec_tlu_pmu_fw_halted;
	assign perfcnt_during_sleep[3:0] = {4 {~(dec_tlu_dbg_halted & dcsr[DCSR_STOPC])}} & {mhpme_vec[39], mhpme_vec[29], mhpme_vec[19], mhpme_vec[9]};
	assign dec_tlu_perfcnt0 = mhpmc_inc_r_d1[0] & ~(perfcnt_halted_d1 & ~perfcnt_during_sleep[0]);
	assign dec_tlu_perfcnt1 = mhpmc_inc_r_d1[1] & ~(perfcnt_halted_d1 & ~perfcnt_during_sleep[1]);
	assign dec_tlu_perfcnt2 = mhpmc_inc_r_d1[2] & ~(perfcnt_halted_d1 & ~perfcnt_during_sleep[2]);
	assign dec_tlu_perfcnt3 = mhpmc_inc_r_d1[3] & ~(perfcnt_halted_d1 & ~perfcnt_during_sleep[3]);
	localparam MHPMC3 = 12'hb03;
	localparam MHPMC3H = 12'hb83;
	assign mhpmc3_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC3);
	assign mhpmc3_wr_en1 = (~perfcnt_halted | perfcnt_during_sleep[0]) & |mhpmc_inc_r[0];
	assign mhpmc3_wr_en = mhpmc3_wr_en0 | mhpmc3_wr_en1;
	assign mhpmc3_incr[63:0] = {mhpmc3h[31:0], mhpmc3[31:0]} + 64'b0000000000000000000000000000000000000000000000000000000000000001;
	assign mhpmc3_ns[31:0] = (mhpmc3_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc3_incr[31:0]);
	rvdffe #(.WIDTH(32)) mhpmc3_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc3_wr_en),
		.din(mhpmc3_ns[31:0]),
		.dout(mhpmc3[31:0])
	);
	assign mhpmc3h_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC3H);
	assign mhpmc3h_wr_en = mhpmc3h_wr_en0 | mhpmc3_wr_en1;
	assign mhpmc3h_ns[31:0] = (mhpmc3h_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc3_incr[63:32]);
	rvdffe #(.WIDTH(32)) mhpmc3h_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc3h_wr_en),
		.din(mhpmc3h_ns[31:0]),
		.dout(mhpmc3h[31:0])
	);
	localparam MHPMC4 = 12'hb04;
	localparam MHPMC4H = 12'hb84;
	assign mhpmc4_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC4);
	assign mhpmc4_wr_en1 = (~perfcnt_halted | perfcnt_during_sleep[1]) & |mhpmc_inc_r[1];
	assign mhpmc4_wr_en = mhpmc4_wr_en0 | mhpmc4_wr_en1;
	assign mhpmc4_incr[63:0] = {mhpmc4h[31:0], mhpmc4[31:0]} + 64'b0000000000000000000000000000000000000000000000000000000000000001;
	assign mhpmc4_ns[31:0] = (mhpmc4_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc4_incr[31:0]);
	rvdffe #(.WIDTH(32)) mhpmc4_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc4_wr_en),
		.din(mhpmc4_ns[31:0]),
		.dout(mhpmc4[31:0])
	);
	assign mhpmc4h_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC4H);
	assign mhpmc4h_wr_en = mhpmc4h_wr_en0 | mhpmc4_wr_en1;
	assign mhpmc4h_ns[31:0] = (mhpmc4h_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc4_incr[63:32]);
	rvdffe #(.WIDTH(32)) mhpmc4h_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc4h_wr_en),
		.din(mhpmc4h_ns[31:0]),
		.dout(mhpmc4h[31:0])
	);
	localparam MHPMC5 = 12'hb05;
	localparam MHPMC5H = 12'hb85;
	assign mhpmc5_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC5);
	assign mhpmc5_wr_en1 = (~perfcnt_halted | perfcnt_during_sleep[2]) & |mhpmc_inc_r[2];
	assign mhpmc5_wr_en = mhpmc5_wr_en0 | mhpmc5_wr_en1;
	assign mhpmc5_incr[63:0] = {mhpmc5h[31:0], mhpmc5[31:0]} + 64'b0000000000000000000000000000000000000000000000000000000000000001;
	assign mhpmc5_ns[31:0] = (mhpmc5_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc5_incr[31:0]);
	rvdffe #(.WIDTH(32)) mhpmc5_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc5_wr_en),
		.din(mhpmc5_ns[31:0]),
		.dout(mhpmc5[31:0])
	);
	assign mhpmc5h_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC5H);
	assign mhpmc5h_wr_en = mhpmc5h_wr_en0 | mhpmc5_wr_en1;
	assign mhpmc5h_ns[31:0] = (mhpmc5h_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc5_incr[63:32]);
	rvdffe #(.WIDTH(32)) mhpmc5h_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc5h_wr_en),
		.din(mhpmc5h_ns[31:0]),
		.dout(mhpmc5h[31:0])
	);
	localparam MHPMC6 = 12'hb06;
	localparam MHPMC6H = 12'hb86;
	assign mhpmc6_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC6);
	assign mhpmc6_wr_en1 = (~perfcnt_halted | perfcnt_during_sleep[3]) & |mhpmc_inc_r[3];
	assign mhpmc6_wr_en = mhpmc6_wr_en0 | mhpmc6_wr_en1;
	assign mhpmc6_incr[63:0] = {mhpmc6h[31:0], mhpmc6[31:0]} + 64'b0000000000000000000000000000000000000000000000000000000000000001;
	assign mhpmc6_ns[31:0] = (mhpmc6_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc6_incr[31:0]);
	rvdffe #(.WIDTH(32)) mhpmc6_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc6_wr_en),
		.din(mhpmc6_ns[31:0]),
		.dout(mhpmc6[31:0])
	);
	assign mhpmc6h_wr_en0 = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPMC6H);
	assign mhpmc6h_wr_en = mhpmc6h_wr_en0 | mhpmc6_wr_en1;
	assign mhpmc6h_ns[31:0] = (mhpmc6h_wr_en0 ? dec_csr_wrdata_r[31:0] : mhpmc6_incr[63:32]);
	rvdffe #(.WIDTH(32)) mhpmc6h_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en(mhpmc6h_wr_en),
		.din(mhpmc6h_ns[31:0]),
		.dout(mhpmc6h[31:0])
	);
	localparam MHPME3 = 12'h323;
	assign zero_event_r = (((((dec_csr_wrdata_r[9:0] > 10'd516) | |dec_csr_wrdata_r[31:10]) | ((dec_csr_wrdata_r[9:0] < 10'd512) & (dec_csr_wrdata_r[9:0] > 10'd56))) | ((dec_csr_wrdata_r[9:0] < 10'd54) & (dec_csr_wrdata_r[9:0] > 10'd50))) | (dec_csr_wrdata_r[9:0] == 10'd29)) | (dec_csr_wrdata_r[9:0] == 10'd33);
	assign event_r[9:0] = (zero_event_r ? {10 {1'sb0}} : dec_csr_wrdata_r[9:0]);
	assign wr_mhpme3_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPME3);
	rvdffe #(.WIDTH(10)) mhpme3_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mhpme3_r),
		.din(event_r[9:0]),
		.dout(mhpme3[9:0])
	);
	localparam MHPME4 = 12'h324;
	assign wr_mhpme4_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPME4);
	rvdffe #(.WIDTH(10)) mhpme4_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mhpme4_r),
		.din(event_r[9:0]),
		.dout(mhpme4[9:0])
	);
	localparam MHPME5 = 12'h325;
	assign wr_mhpme5_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPME5);
	rvdffe #(.WIDTH(10)) mhpme5_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mhpme5_r),
		.din(event_r[9:0]),
		.dout(mhpme5[9:0])
	);
	localparam MHPME6 = 12'h326;
	assign wr_mhpme6_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MHPME6);
	rvdffe #(.WIDTH(10)) mhpme6_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mhpme6_r),
		.din(event_r[9:0]),
		.dout(mhpme6[9:0])
	);
	localparam MCOUNTINHIBIT = 12'h320;
	assign wr_mcountinhibit_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MCOUNTINHIBIT);
	rvdffs #(.WIDTH(6)) mcountinhibit_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.en(wr_mcountinhibit_r),
		.din({dec_csr_wrdata_r[6:2], dec_csr_wrdata_r[0]}),
		.dout({mcountinhibit[6:2], mcountinhibit[0]})
	);
	assign mcountinhibit[1] = 1'b0;
	wire [4:0] dec_tlu_exc_cause_wb1_raw;
	wire [4:0] dec_tlu_exc_cause_wb2;
	wire dec_tlu_int_valid_wb1_raw;
	wire dec_tlu_int_valid_wb2;
	assign {dec_tlu_i0_valid_wb1, dec_tlu_i0_exc_valid_wb1, dec_tlu_exc_cause_wb1_raw[4:0], dec_tlu_int_valid_wb1_raw} = {8 {~dec_tlu_trace_disable}} & {i0_valid_wb, (i0_exception_valid_r_d1 | lsu_i0_exc_r_d1) | (trigger_hit_r_d1 & ~trigger_hit_dmode_r_d1), exc_cause_wb[4:0], interrupt_valid_r_d1};
	rvdffie #(
		.WIDTH(6),
		.OVERRIDE(1)
	) traceskidff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din({dec_tlu_exc_cause_wb1_raw[4:0], dec_tlu_int_valid_wb1_raw}),
		.dout({dec_tlu_exc_cause_wb2[4:0], dec_tlu_int_valid_wb2})
	);
	assign dec_tlu_exc_cause_wb1[4:0] = (dec_tlu_int_valid_wb2 ? dec_tlu_exc_cause_wb2[4:0] : dec_tlu_exc_cause_wb1_raw[4:0]);
	assign dec_tlu_int_valid_wb1 = dec_tlu_int_valid_wb2;
	assign dec_tlu_mtval_wb1 = mtval[31:0];
	assign csr_misa = (((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_mvendorid = ((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_marchid = ((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mimpid = ((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mhartid = (dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[2];
	assign csr_mstatus = (((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0];
	assign csr_mtvec = (((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_mip = (!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[2];
	assign csr_mie = (((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0];
	assign csr_mcyclel = ((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1];
	assign csr_mcycleh = (((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1];
	assign csr_minstretl = (((((!dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_minstreth = (((((!dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mscratch = (((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mepc = ((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mcause = ((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mscause = (dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2];
	assign csr_mtval = ((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mrac = ((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1];
	assign csr_dmst = (((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1];
	assign csr_mdseac = ((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3];
	assign csr_meihap = (dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[3];
	assign csr_meivt = ((((!dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_meipt = ((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_meicurpl = (dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[2];
	assign csr_meicidpl = ((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_dcsr = (((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[0];
	assign csr_mcgc = ((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[0];
	assign csr_mfdc = (((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_dpc = (((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[0];
	assign csr_mtsel = (((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mtdata1 = ((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[0];
	assign csr_mtdata2 = ((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[1];
	assign csr_mhpmc3 = ((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_mhpmc4 = (((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mhpmc5 = ((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mhpmc6 = (((((!dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mhpmc3h = ((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mhpmc4h = (((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mhpmc5h = ((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mhpmc6h = (((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mhpme3 = ((((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_mhpme4 = ((((dec_csr_rdaddr_d[5] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mhpme5 = ((((dec_csr_rdaddr_d[5] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mhpme6 = ((((dec_csr_rdaddr_d[5] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mcountinhibit = ((((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0];
	assign csr_mitctl0 = (((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mitctl1 = (((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mitb0 = (((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_mitb1 = (((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mitcnt0 = (((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0];
	assign csr_mitcnt1 = ((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_mpmc = (((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1];
	assign csr_meicpct = ((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_micect = (((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_miccmect = ((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[0];
	assign csr_mdccmect = ((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mfdht = (((dec_csr_rdaddr_d[6] & dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_mfdhs = ((dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0];
	assign csr_dicawics = ((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_dicad0h = ((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1];
	assign csr_dicad0 = (((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign csr_dicad1 = (((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0];
	assign csr_dicago = (((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0];
	assign presync = ((((((((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0]) | (((((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0])) | (((((!dec_csr_rdaddr_d[6] & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1])) | ((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1])) | ((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | (((((dec_csr_rdaddr_d[7] & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]);
	assign postsync = (((((((((dec_csr_rdaddr_d[10] & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0]) | ((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0])) | (((!dec_csr_rdaddr_d[7] & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0])) | (((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[0])) | ((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0])) | (((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1])) | ((((dec_csr_rdaddr_d[10] & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]);
	assign legal = (((((((((((((((((((((((((((((((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0]) | (((((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1])) | ((((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | (((((((((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | ((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[0])) | (((((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1])) | (((((((((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[0])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1])) | (((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2])) | ((((((((((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[1])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[2])) | (((((((((dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & dec_csr_rdaddr_d[1])) | ((((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[1]) & dec_csr_rdaddr_d[0])) | ((((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2])) | (((((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | ((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[2])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & dec_csr_rdaddr_d[1])) | ((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[0])) | (((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2])) | ((((((((((!dec_csr_rdaddr_d[11] & dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2]) & !dec_csr_rdaddr_d[0])) | ((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[1])) | (((((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[2])) | (((((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[5]) & !dec_csr_rdaddr_d[4]) & !dec_csr_rdaddr_d[3]) & !dec_csr_rdaddr_d[1]) & !dec_csr_rdaddr_d[0])) | (((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[3])) | ((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[3])) | (((((((!dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[7]) & !dec_csr_rdaddr_d[6]) & dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4])) | ((((((dec_csr_rdaddr_d[11] & !dec_csr_rdaddr_d[10]) & dec_csr_rdaddr_d[9]) & dec_csr_rdaddr_d[8]) & !dec_csr_rdaddr_d[6]) & !dec_csr_rdaddr_d[5]) & dec_csr_rdaddr_d[4]);
	assign dec_tlu_presync_d = (presync & dec_csr_any_unq_d) & ~dec_csr_wen_unq_d;
	assign dec_tlu_postsync_d = postsync & dec_csr_any_unq_d;
	assign conditionally_illegal = (((((csr_mitcnt0 | csr_mitcnt1) | csr_mitb0) | csr_mitb1) | csr_mitctl0) | csr_mitctl1) & !pt[4-:5];
	assign valid_csr = ((legal & (~(((((((csr_dcsr | csr_dpc) | csr_dmst) | csr_dicawics) | csr_dicad0) | csr_dicad0h) | csr_dicad1) | csr_dicago) | dbg_tlu_halted_f)) & ~fast_int_meicpct) & ~conditionally_illegal;
	assign dec_csr_legal_d = (dec_csr_any_unq_d & valid_csr) & ~(dec_csr_wen_unq_d & (((((csr_mvendorid | csr_marchid) | csr_mimpid) | csr_mhartid) | csr_mdseac) | csr_meihap));
	assign dec_csr_rddata_d[31:0] = ((((((((((((((((((((((((((((((((((((((((((((((((((((((({32 {csr_misa}} & 32'h40201104) | ({32 {csr_mvendorid}} & 32'h00000045)) | ({32 {csr_marchid}} & 32'h00000010)) | ({32 {csr_mimpid}} & 32'h00000003)) | ({32 {csr_mhartid}} & {core_id[31:4], 4'b0000})) | ({32 {csr_mstatus}} & {{15 {1'b0}}, 2'b01, 2'b00, 2'b11, 3'b000, mstatus[1], 3'b000, mstatus[0], 3'b000})) | ({32 {csr_mtvec}} & {mtvec[30:1], 1'b0, mtvec[0]})) | ({32 {csr_mip}} & {1'b0, mip[5:3], 16'b0000000000000000, mip[2], 3'b000, mip[1], 3'b000, mip[0], 3'b000})) | ({32 {csr_mie}} & {1'b0, mie[5:3], 16'b0000000000000000, mie[2], 3'b000, mie[1], 3'b000, mie[0], 3'b000})) | ({32 {csr_mcyclel}} & mcyclel[31:0])) | ({32 {csr_mcycleh}} & mcycleh_inc[31:0])) | ({32 {csr_minstretl}} & minstretl_read[31:0])) | ({32 {csr_minstreth}} & minstreth_read[31:0])) | ({32 {csr_mscratch}} & mscratch[31:0])) | ({32 {csr_mepc}} & {mepc[31:1], 1'b0})) | ({32 {csr_mcause}} & mcause[31:0])) | ({32 {csr_mscause}} & {28'b0000000000000000000000000000, mscause[3:0]})) | ({32 {csr_mtval}} & mtval[31:0])) | ({32 {csr_mrac}} & mrac[31:0])) | ({32 {csr_mdseac}} & mdseac[31:0])) | ({32 {csr_meivt}} & {meivt[31:10], 10'b0000000000})) | ({32 {csr_meihap}} & {meivt[31:10], meihap[9:2], 2'b00})) | ({32 {csr_meicurpl}} & {28'b0000000000000000000000000000, meicurpl[3:0]})) | ({32 {csr_meicidpl}} & {28'b0000000000000000000000000000, meicidpl[3:0]})) | ({32 {csr_meipt}} & {28'b0000000000000000000000000000, meipt[3:0]})) | ({32 {csr_mcgc}} & {22'b0000000000000000000000, mcgc[9:0]})) | ({32 {csr_mfdc}} & {13'b0000000000000, mfdc[18:0]})) | ({32 {csr_dcsr}} & {16'h4000, dcsr[15:2], 2'b11})) | ({32 {csr_dpc}} & {dpc[31:1], 1'b0})) | ({32 {csr_dicad0}} & dicad0[31:0])) | ({32 {csr_dicad0h}} & dicad0h[31:0])) | ({32 {csr_dicad1}} & dicad1[31:0])) | ({32 {csr_dicawics}} & {7'b0000000, dicawics[16], 2'b00, dicawics[15:14], 3'b000, dicawics[13:0], 3'b000})) | ({32 {csr_mtsel}} & {30'b000000000000000000000000000000, mtsel[1:0]})) | ({32 {csr_mtdata1}} & {mtdata1_tsel_out[31:0]})) | ({32 {csr_mtdata2}} & {mtdata2_tsel_out[31:0]})) | ({32 {csr_micect}} & {micect[31:0]})) | ({32 {csr_miccmect}} & {miccmect[31:0]})) | ({32 {csr_mdccmect}} & {mdccmect[31:0]})) | ({32 {csr_mhpmc3}} & mhpmc3[31:0])) | ({32 {csr_mhpmc4}} & mhpmc4[31:0])) | ({32 {csr_mhpmc5}} & mhpmc5[31:0])) | ({32 {csr_mhpmc6}} & mhpmc6[31:0])) | ({32 {csr_mhpmc3h}} & mhpmc3h[31:0])) | ({32 {csr_mhpmc4h}} & mhpmc4h[31:0])) | ({32 {csr_mhpmc5h}} & mhpmc5h[31:0])) | ({32 {csr_mhpmc6h}} & mhpmc6h[31:0])) | ({32 {csr_mfdht}} & {26'b00000000000000000000000000, mfdht[5:0]})) | ({32 {csr_mfdhs}} & {30'b000000000000000000000000000000, mfdhs[1:0]})) | ({32 {csr_mhpme3}} & {22'b0000000000000000000000, mhpme3[9:0]})) | ({32 {csr_mhpme4}} & {22'b0000000000000000000000, mhpme4[9:0]})) | ({32 {csr_mhpme5}} & {22'b0000000000000000000000, mhpme5[9:0]})) | ({32 {csr_mhpme6}} & {22'b0000000000000000000000, mhpme6[9:0]})) | ({32 {csr_mcountinhibit}} & {25'b0000000000000000000000000, mcountinhibit[6:0]})) | ({32 {csr_mpmc}} & {30'b000000000000000000000000000000, mpmc[1], 1'b0})) | ({32 {dec_timer_read_d}} & dec_timer_rddata_d[31:0]);
endmodule
module eb1_dec_timer_ctl (
	clk,
	free_l2clk,
	csr_wr_clk,
	rst_l,
	dec_csr_wen_r_mod,
	dec_csr_wraddr_r,
	dec_csr_wrdata_r,
	csr_mitctl0,
	csr_mitctl1,
	csr_mitb0,
	csr_mitb1,
	csr_mitcnt0,
	csr_mitcnt1,
	dec_pause_state,
	dec_tlu_pmu_fw_halted,
	internal_dbg_halt_timers,
	dec_timer_rddata_d,
	dec_timer_read_d,
	dec_timer_t0_pulse,
	dec_timer_t1_pulse,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire free_l2clk;
	input wire csr_wr_clk;
	input wire rst_l;
	input wire dec_csr_wen_r_mod;
	input wire [11:0] dec_csr_wraddr_r;
	input wire [31:0] dec_csr_wrdata_r;
	input wire csr_mitctl0;
	input wire csr_mitctl1;
	input wire csr_mitb0;
	input wire csr_mitb1;
	input wire csr_mitcnt0;
	input wire csr_mitcnt1;
	input wire dec_pause_state;
	input wire dec_tlu_pmu_fw_halted;
	input wire internal_dbg_halt_timers;
	output wire [31:0] dec_timer_rddata_d;
	output wire dec_timer_read_d;
	output wire dec_timer_t0_pulse;
	output wire dec_timer_t1_pulse;
	input wire scan_mode;
	localparam MITCTL_ENABLE = 0;
	localparam MITCTL_ENABLE_HALTED = 1;
	localparam MITCTL_ENABLE_PAUSED = 2;
	wire [31:0] mitcnt0_ns;
	wire [31:0] mitcnt0;
	wire [31:0] mitcnt1_ns;
	wire [31:0] mitcnt1;
	wire [31:0] mitb0;
	wire [31:0] mitb1;
	wire [31:0] mitb0_b;
	wire [31:0] mitb1_b;
	wire [31:0] mitcnt0_inc;
	wire [31:0] mitcnt1_inc;
	wire [2:0] mitctl0_ns;
	wire [2:0] mitctl0;
	wire [3:0] mitctl1_ns;
	wire [3:0] mitctl1;
	wire wr_mitcnt0_r;
	wire wr_mitcnt1_r;
	wire wr_mitb0_r;
	wire wr_mitb1_r;
	wire wr_mitctl0_r;
	wire wr_mitctl1_r;
	wire mitcnt0_inc_ok;
	wire mitcnt1_inc_ok;
	wire mitcnt0_inc_cout;
	wire mitcnt1_inc_cout;
	wire mit0_match_ns;
	wire mit1_match_ns;
	wire mitctl0_0_b_ns;
	wire mitctl0_0_b;
	wire mitctl1_0_b_ns;
	wire mitctl1_0_b;
	assign mit0_match_ns = mitcnt0[31:0] >= mitb0[31:0];
	assign mit1_match_ns = mitcnt1[31:0] >= mitb1[31:0];
	assign dec_timer_t0_pulse = mit0_match_ns;
	assign dec_timer_t1_pulse = mit1_match_ns;
	localparam MITCNT0 = 12'h7d2;
	assign wr_mitcnt0_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITCNT0);
	assign mitcnt0_inc_ok = ((mitctl0[MITCTL_ENABLE] & (~dec_pause_state | mitctl0[MITCTL_ENABLE_PAUSED])) & (~dec_tlu_pmu_fw_halted | mitctl0[MITCTL_ENABLE_HALTED])) & ~internal_dbg_halt_timers;
	assign {mitcnt0_inc_cout, mitcnt0_inc[7:0]} = mitcnt0[7:0] + 8'b00000001;
	assign mitcnt0_inc[31:8] = mitcnt0[31:8] + {23'b00000000000000000000000, mitcnt0_inc_cout};
	assign mitcnt0_ns[31:0] = (wr_mitcnt0_r ? dec_csr_wrdata_r[31:0] : (mit0_match_ns ? 'b0 : mitcnt0_inc[31:0]));
	rvdffe #(.WIDTH(24)) mitcnt0_ffb(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en((wr_mitcnt0_r | (mitcnt0_inc_ok & mitcnt0_inc_cout)) | mit0_match_ns),
		.din(mitcnt0_ns[31:8]),
		.dout(mitcnt0[31:8])
	);
	rvdffe #(.WIDTH(8)) mitcnt0_ffa(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en((wr_mitcnt0_r | mitcnt0_inc_ok) | mit0_match_ns),
		.din(mitcnt0_ns[7:0]),
		.dout(mitcnt0[7:0])
	);
	localparam MITCNT1 = 12'h7d5;
	assign wr_mitcnt1_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITCNT1);
	assign mitcnt1_inc_ok = (((mitctl1[MITCTL_ENABLE] & (~dec_pause_state | mitctl1[MITCTL_ENABLE_PAUSED])) & (~dec_tlu_pmu_fw_halted | mitctl1[MITCTL_ENABLE_HALTED])) & ~internal_dbg_halt_timers) & (~mitctl1[3] | mit0_match_ns);
	assign {mitcnt1_inc_cout, mitcnt1_inc[7:0]} = mitcnt1[7:0] + 8'b00000001;
	assign mitcnt1_inc[31:8] = mitcnt1[31:8] + {23'b00000000000000000000000, mitcnt1_inc_cout};
	assign mitcnt1_ns[31:0] = (wr_mitcnt1_r ? dec_csr_wrdata_r[31:0] : (mit1_match_ns ? 'b0 : mitcnt1_inc[31:0]));
	rvdffe #(.WIDTH(24)) mitcnt1_ffb(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en((wr_mitcnt1_r | (mitcnt1_inc_ok & mitcnt1_inc_cout)) | mit1_match_ns),
		.din(mitcnt1_ns[31:8]),
		.dout(mitcnt1[31:8])
	);
	rvdffe #(.WIDTH(8)) mitcnt1_ffa(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.en((wr_mitcnt1_r | mitcnt1_inc_ok) | mit1_match_ns),
		.din(mitcnt1_ns[7:0]),
		.dout(mitcnt1[7:0])
	);
	localparam MITB0 = 12'h7d3;
	assign wr_mitb0_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITB0);
	rvdffe #(.WIDTH(32)) mitb0_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mitb0_r),
		.din(~dec_csr_wrdata_r[31:0]),
		.dout(mitb0_b[31:0])
	);
	assign mitb0[31:0] = ~mitb0_b[31:0];
	localparam MITB1 = 12'h7d6;
	assign wr_mitb1_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITB1);
	rvdffe #(.WIDTH(32)) mitb1_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(wr_mitb1_r),
		.din(~dec_csr_wrdata_r[31:0]),
		.dout(mitb1_b[31:0])
	);
	assign mitb1[31:0] = ~mitb1_b[31:0];
	localparam MITCTL0 = 12'h7d4;
	assign wr_mitctl0_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITCTL0);
	assign mitctl0_ns[2:0] = (wr_mitctl0_r ? {dec_csr_wrdata_r[2:0]} : {mitctl0[2:0]});
	assign mitctl0_0_b_ns = ~mitctl0_ns[0];
	rvdffs #(.WIDTH(3)) mitctl0_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.en(wr_mitctl0_r),
		.din({mitctl0_ns[2:1], mitctl0_0_b_ns}),
		.dout({mitctl0[2:1], mitctl0_0_b})
	);
	assign mitctl0[0] = ~mitctl0_0_b;
	localparam MITCTL1 = 12'h7d7;
	assign wr_mitctl1_r = dec_csr_wen_r_mod & (dec_csr_wraddr_r[11:0] == MITCTL1);
	assign mitctl1_ns[3:0] = (wr_mitctl1_r ? {dec_csr_wrdata_r[3:0]} : {mitctl1[3:0]});
	assign mitctl1_0_b_ns = ~mitctl1_ns[0];
	rvdffs #(.WIDTH(4)) mitctl1_ff(
		.rst_l(rst_l),
		.clk(csr_wr_clk),
		.en(wr_mitctl1_r),
		.din({mitctl1_ns[3:1], mitctl1_0_b_ns}),
		.dout({mitctl1[3:1], mitctl1_0_b})
	);
	assign mitctl1[0] = ~mitctl1_0_b;
	assign dec_timer_read_d = ((((csr_mitcnt1 | csr_mitcnt0) | csr_mitb1) | csr_mitb0) | csr_mitctl0) | csr_mitctl1;
	assign dec_timer_rddata_d[31:0] = ((((({32 {csr_mitcnt0}} & mitcnt0[31:0]) | ({32 {csr_mitcnt1}} & mitcnt1[31:0])) | ({32 {csr_mitb0}} & mitb0[31:0])) | ({32 {csr_mitb1}} & mitb1[31:0])) | ({32 {csr_mitctl0}} & {29'b00000000000000000000000000000, mitctl0[2:0]})) | ({32 {csr_mitctl1}} & {28'b0000000000000000000000000000, mitctl1[3:0]});
endmodule
module eb1_dec_trigger (
	trigger_pkt_any,
	dec_i0_pc_d,
	dec_i0_trigger_match_d
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [151:0] trigger_pkt_any;
	input wire [31:1] dec_i0_pc_d;
	output wire [3:0] dec_i0_trigger_match_d;
	wire [127:0] dec_i0_match_data;
	wire [3:0] dec_i0_trigger_data_match;
	generate
		genvar i;
		for (i = 0; i < 4; i = i + 1) begin
			assign dec_i0_match_data[(i * 32) + 31-:32] = {32 {~trigger_pkt_any[(i * 38) + 37] & trigger_pkt_any[(i * 38) + 33]}} & {dec_i0_pc_d[31:1], trigger_pkt_any[i * 38]};
			rvmaskandmatch trigger_i0_match(
				.mask(trigger_pkt_any[(i * 38) + 31-:32]),
				.data(dec_i0_match_data[(i * 32) + 31-:32]),
				.masken(trigger_pkt_any[(i * 38) + 36]),
				.match(dec_i0_trigger_data_match[i])
			);
			assign dec_i0_trigger_match_d[i] = (trigger_pkt_any[(i * 38) + 33] & trigger_pkt_any[(i * 38) + 32]) & dec_i0_trigger_data_match[i];
		end
	endgenerate
endmodule
module eb1_exu (
	clk,
	rst_l,
	scan_mode,
	dec_data_en,
	dec_ctl_en,
	dbg_cmd_wrdata,
	i0_ap,
	dec_debug_wdata_rs1_d,
	dec_i0_predict_p_d,
	i0_predict_fghr_d,
	i0_predict_index_d,
	i0_predict_btag_d,
	lsu_result_m,
	lsu_nonblock_load_data,
	dec_i0_rs1_en_d,
	dec_i0_rs2_en_d,
	gpr_i0_rs1_d,
	gpr_i0_rs2_d,
	dec_i0_immed_d,
	dec_i0_result_r,
	dec_i0_br_immed_d,
	dec_i0_alu_decode_d,
	dec_i0_branch_d,
	dec_i0_select_pc_d,
	dec_i0_pc_d,
	dec_i0_rs1_bypass_en_d,
	dec_i0_rs2_bypass_en_d,
	dec_csr_ren_d,
	dec_csr_rddata_d,
	dec_qual_lsu_d,
	mul_p,
	div_p,
	dec_div_cancel,
	pred_correct_npc_x,
	dec_tlu_flush_lower_r,
	dec_tlu_flush_path_r,
	dec_extint_stall,
	dec_tlu_meihap,
	exu_lsu_rs1_d,
	exu_lsu_rs2_d,
	exu_flush_final,
	exu_flush_path_final,
	exu_i0_result_x,
	exu_i0_pc_x,
	exu_csr_rs1_x,
	exu_npc_r,
	exu_i0_br_hist_r,
	exu_i0_br_error_r,
	exu_i0_br_start_error_r,
	exu_i0_br_index_r,
	exu_i0_br_valid_r,
	exu_i0_br_mp_r,
	exu_i0_br_middle_r,
	exu_i0_br_fghr_r,
	exu_i0_br_way_r,
	exu_mp_pkt,
	exu_mp_eghr,
	exu_mp_fghr,
	exu_mp_index,
	exu_mp_btag,
	exu_pmu_i0_br_misp,
	exu_pmu_i0_br_ataken,
	exu_pmu_i0_pc4,
	exu_div_result,
	exu_div_wren
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire [1:0] dec_data_en;
	input wire [1:0] dec_ctl_en;
	input wire [31:0] dbg_cmd_wrdata;
	input wire [43:0] i0_ap;
	input wire dec_debug_wdata_rs1_d;
	input wire [55:0] dec_i0_predict_p_d;
	input wire [pt[2236-:8] - 1:0] i0_predict_fghr_d;
	input wire [pt[2172-:9]:pt[2163-:6]] i0_predict_index_d;
	input wire [pt[2139-:9] - 1:0] i0_predict_btag_d;
	input wire [31:0] lsu_result_m;
	input wire [31:0] lsu_nonblock_load_data;
	input wire dec_i0_rs1_en_d;
	input wire dec_i0_rs2_en_d;
	input wire [31:0] gpr_i0_rs1_d;
	input wire [31:0] gpr_i0_rs2_d;
	input wire [31:0] dec_i0_immed_d;
	input wire [31:0] dec_i0_result_r;
	input wire [12:1] dec_i0_br_immed_d;
	input wire dec_i0_alu_decode_d;
	input wire dec_i0_branch_d;
	input wire dec_i0_select_pc_d;
	input wire [31:1] dec_i0_pc_d;
	input wire [3:0] dec_i0_rs1_bypass_en_d;
	input wire [3:0] dec_i0_rs2_bypass_en_d;
	input wire dec_csr_ren_d;
	input wire [31:0] dec_csr_rddata_d;
	input wire dec_qual_lsu_d;
	input wire [19:0] mul_p;
	input wire [2:0] div_p;
	input wire dec_div_cancel;
	input wire [31:1] pred_correct_npc_x;
	input wire dec_tlu_flush_lower_r;
	input wire [31:1] dec_tlu_flush_path_r;
	input wire dec_extint_stall;
	input wire [31:2] dec_tlu_meihap;
	output wire [31:0] exu_lsu_rs1_d;
	output wire [31:0] exu_lsu_rs2_d;
	output wire exu_flush_final;
	output wire [31:1] exu_flush_path_final;
	output wire [31:0] exu_i0_result_x;
	output wire [31:1] exu_i0_pc_x;
	output wire [31:0] exu_csr_rs1_x;
	output wire [31:1] exu_npc_r;
	output wire [1:0] exu_i0_br_hist_r;
	output wire exu_i0_br_error_r;
	output wire exu_i0_br_start_error_r;
	output wire [pt[2172-:9]:pt[2163-:6]] exu_i0_br_index_r;
	output wire exu_i0_br_valid_r;
	output wire exu_i0_br_mp_r;
	output wire exu_i0_br_middle_r;
	output wire [pt[2236-:8] - 1:0] exu_i0_br_fghr_r;
	output wire exu_i0_br_way_r;
	output wire [55:0] exu_mp_pkt;
	output wire [pt[2236-:8] - 1:0] exu_mp_eghr;
	output wire [pt[2236-:8] - 1:0] exu_mp_fghr;
	output wire [pt[2172-:9]:pt[2163-:6]] exu_mp_index;
	output wire [pt[2139-:9] - 1:0] exu_mp_btag;
	output wire exu_pmu_i0_br_misp;
	output wire exu_pmu_i0_br_ataken;
	output wire exu_pmu_i0_pc4;
	output wire [31:0] exu_div_result;
	output wire exu_div_wren;
	wire [31:0] i0_rs1_bypass_data_d;
	wire [31:0] i0_rs2_bypass_data_d;
	wire i0_rs1_bypass_en_d;
	wire i0_rs2_bypass_en_d;
	wire [31:0] i0_rs1_d;
	wire [31:0] i0_rs2_d;
	wire [31:0] muldiv_rs1_d;
	wire [31:1] pred_correct_npc_r;
	wire i0_pred_correct_upper_r;
	wire [31:1] i0_flush_path_upper_r;
	wire x_data_en;
	wire x_data_en_q1;
	wire x_data_en_q2;
	wire r_data_en;
	wire r_data_en_q2;
	wire x_ctl_en;
	wire r_ctl_en;
	wire [pt[2236-:8] - 1:0] ghr_d_ns;
	wire [pt[2236-:8] - 1:0] ghr_d;
	wire [pt[2236-:8] - 1:0] ghr_x_ns;
	wire [pt[2236-:8] - 1:0] ghr_x;
	wire i0_taken_d;
	wire i0_taken_x;
	wire i0_valid_d;
	wire i0_valid_x;
	wire [pt[2236-:8] - 1:0] after_flush_eghr;
	wire [55:0] final_predict_mp;
	reg [55:0] i0_predict_newp_d;
	wire flush_in_d;
	wire [31:0] alu_result_x;
	wire mul_valid_x;
	wire [31:0] mul_result_x;
	wire [55:0] i0_pp_r;
	wire i0_flush_upper_d;
	wire [31:1] i0_flush_path_d;
	wire [55:0] i0_predict_p_d;
	wire i0_pred_correct_upper_d;
	wire i0_flush_upper_x;
	wire [31:1] i0_flush_path_x;
	wire [55:0] i0_predict_p_x;
	wire i0_pred_correct_upper_x;
	wire i0_branch_x;
	localparam PREDPIPESIZE = (((pt[2172-:9] - pt[2163-:6]) + 1) + pt[2236-:8]) + pt[2139-:9];
	wire [PREDPIPESIZE - 1:0] predpipe_d;
	wire [PREDPIPESIZE - 1:0] predpipe_x;
	wire [PREDPIPESIZE - 1:0] predpipe_r;
	wire [PREDPIPESIZE - 1:0] final_predpipe_mp;
	rvdffpcie #(.WIDTH(31)) i_flush_path_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(x_data_en),
		.din(i0_flush_path_d[31:1]),
		.dout(i0_flush_path_x[31:1])
	);
	rvdffe #(.WIDTH(32)) i_csr_rs1_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(x_data_en_q1),
		.din(i0_rs1_d[31:0]),
		.dout(exu_csr_rs1_x[31:0])
	);
	rvdffppe #(.WIDTH(56)) i_predictpacket_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(x_data_en),
		.din(i0_predict_p_d),
		.dout(i0_predict_p_x)
	);
	rvdffe #(.WIDTH(PREDPIPESIZE)) i_predpipe_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(x_data_en_q2),
		.din(predpipe_d),
		.dout(predpipe_x)
	);
	rvdffe #(.WIDTH(PREDPIPESIZE)) i_predpipe_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(r_data_en_q2),
		.din(predpipe_x),
		.dout(predpipe_r)
	);
	rvdffe #(.WIDTH(4 + pt[2236-:8])) i_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(x_ctl_en),
		.din({i0_valid_d, i0_taken_d, i0_flush_upper_d, i0_pred_correct_upper_d, ghr_x_ns[pt[2236-:8] - 1:0]}),
		.dout({i0_valid_x, i0_taken_x, i0_flush_upper_x, i0_pred_correct_upper_x, ghr_x[pt[2236-:8] - 1:0]})
	);
	rvdffppe #(.WIDTH(57)) i_r_ff0(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(r_ctl_en),
		.din({i0_pred_correct_upper_x, i0_predict_p_x}),
		.dout({i0_pred_correct_upper_r, i0_pp_r})
	);
	rvdffpcie #(.WIDTH(31)) i_flush_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(r_data_en),
		.din(i0_flush_path_x[31:1]),
		.dout(i0_flush_path_upper_r[31:1])
	);
	rvdffpcie #(.WIDTH(31)) i_npc_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(r_data_en),
		.din(pred_correct_npc_x[31:1]),
		.dout(pred_correct_npc_r[31:1])
	);
	rvdffie #(
		.WIDTH(pt[2236-:8] + 2),
		.OVERRIDE(1)
	) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din({ghr_d_ns[pt[2236-:8] - 1:0], mul_p[19], dec_i0_branch_d}),
		.dout({ghr_d[pt[2236-:8] - 1:0], mul_valid_x, i0_branch_x})
	);
	assign predpipe_d[PREDPIPESIZE - 1:0] = {i0_predict_fghr_d, i0_predict_index_d, i0_predict_btag_d};
	assign i0_rs1_bypass_en_d = ((dec_i0_rs1_bypass_en_d[0] | dec_i0_rs1_bypass_en_d[1]) | dec_i0_rs1_bypass_en_d[2]) | dec_i0_rs1_bypass_en_d[3];
	assign i0_rs2_bypass_en_d = ((dec_i0_rs2_bypass_en_d[0] | dec_i0_rs2_bypass_en_d[1]) | dec_i0_rs2_bypass_en_d[2]) | dec_i0_rs2_bypass_en_d[3];
	assign i0_rs1_bypass_data_d[31:0] = ((({32 {dec_i0_rs1_bypass_en_d[0]}} & dec_i0_result_r[31:0]) | ({32 {dec_i0_rs1_bypass_en_d[1]}} & lsu_result_m[31:0])) | ({32 {dec_i0_rs1_bypass_en_d[2]}} & exu_i0_result_x[31:0])) | ({32 {dec_i0_rs1_bypass_en_d[3]}} & lsu_nonblock_load_data[31:0]);
	assign i0_rs2_bypass_data_d[31:0] = ((({32 {dec_i0_rs2_bypass_en_d[0]}} & dec_i0_result_r[31:0]) | ({32 {dec_i0_rs2_bypass_en_d[1]}} & lsu_result_m[31:0])) | ({32 {dec_i0_rs2_bypass_en_d[2]}} & exu_i0_result_x[31:0])) | ({32 {dec_i0_rs2_bypass_en_d[3]}} & lsu_nonblock_load_data[31:0]);
	assign i0_rs1_d[31:0] = ((({32 {i0_rs1_bypass_en_d}} & i0_rs1_bypass_data_d[31:0]) | ({32 {~i0_rs1_bypass_en_d & dec_i0_select_pc_d}} & {dec_i0_pc_d[31:1], 1'b0})) | ({32 {~i0_rs1_bypass_en_d & dec_debug_wdata_rs1_d}} & dbg_cmd_wrdata[31:0])) | ({32 {(~i0_rs1_bypass_en_d & ~dec_debug_wdata_rs1_d) & dec_i0_rs1_en_d}} & gpr_i0_rs1_d[31:0]);
	assign i0_rs2_d[31:0] = (({32 {~i0_rs2_bypass_en_d & dec_i0_rs2_en_d}} & gpr_i0_rs2_d[31:0]) | ({32 {~i0_rs2_bypass_en_d}} & dec_i0_immed_d[31:0])) | ({32 {i0_rs2_bypass_en_d}} & i0_rs2_bypass_data_d[31:0]);
	assign exu_lsu_rs1_d[31:0] = (({32 {((~i0_rs1_bypass_en_d & ~dec_extint_stall) & dec_i0_rs1_en_d) & dec_qual_lsu_d}} & gpr_i0_rs1_d[31:0]) | ({32 {(i0_rs1_bypass_en_d & ~dec_extint_stall) & dec_qual_lsu_d}} & i0_rs1_bypass_data_d[31:0])) | ({32 {dec_extint_stall & dec_qual_lsu_d}} & {dec_tlu_meihap[31:2], 2'b00});
	assign exu_lsu_rs2_d[31:0] = ({32 {((~i0_rs2_bypass_en_d & ~dec_extint_stall) & dec_i0_rs2_en_d) & dec_qual_lsu_d}} & gpr_i0_rs2_d[31:0]) | ({32 {(i0_rs2_bypass_en_d & ~dec_extint_stall) & dec_qual_lsu_d}} & i0_rs2_bypass_data_d[31:0]);
	assign muldiv_rs1_d[31:0] = ({32 {~i0_rs1_bypass_en_d & dec_i0_rs1_en_d}} & gpr_i0_rs1_d[31:0]) | ({32 {i0_rs1_bypass_en_d}} & i0_rs1_bypass_data_d[31:0]);
	assign x_data_en = dec_data_en[1];
	assign x_data_en_q1 = dec_data_en[1] & dec_csr_ren_d;
	assign x_data_en_q2 = dec_data_en[1] & dec_i0_branch_d;
	assign r_data_en = dec_data_en[0];
	assign r_data_en_q2 = dec_data_en[0] & i0_branch_x;
	assign x_ctl_en = dec_ctl_en[1];
	assign r_ctl_en = dec_ctl_en[0];
	eb1_exu_alu_ctl #(.pt(pt)) i_alu(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.enable(x_data_en),
		.pp_in(i0_predict_newp_d),
		.valid_in(dec_i0_alu_decode_d),
		.flush_upper_x(i0_flush_upper_x),
		.flush_lower_r(dec_tlu_flush_lower_r),
		.a_in(i0_rs1_d[31:0]),
		.b_in(i0_rs2_d[31:0]),
		.pc_in(dec_i0_pc_d[31:1]),
		.brimm_in(dec_i0_br_immed_d[12:1]),
		.ap(i0_ap),
		.csr_ren_in(dec_csr_ren_d),
		.csr_rddata_in(dec_csr_rddata_d[31:0]),
		.result_ff(alu_result_x[31:0]),
		.flush_upper_out(i0_flush_upper_d),
		.flush_final_out(exu_flush_final),
		.flush_path_out(i0_flush_path_d[31:1]),
		.predict_p_out(i0_predict_p_d),
		.pred_correct_out(i0_pred_correct_upper_d),
		.pc_ff(exu_i0_pc_x[31:1])
	);
	eb1_exu_mul_ctl #(.pt(pt)) i_mul(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.mul_p(mul_p & {20 {mul_p[19]}}),
		.rs1_in(muldiv_rs1_d[31:0] & {32 {mul_p[19]}}),
		.rs2_in(i0_rs2_d[31:0] & {32 {mul_p[19]}}),
		.result_x(mul_result_x[31:0])
	);
	eb1_exu_div_ctl #(.pt(pt)) i_div(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.cancel(dec_div_cancel),
		.dp(div_p),
		.dividend(muldiv_rs1_d[31:0]),
		.divisor(i0_rs2_d[31:0]),
		.finish_dly(exu_div_wren),
		.out(exu_div_result[31:0])
	);
	assign exu_i0_result_x[31:0] = (mul_valid_x ? mul_result_x[31:0] : alu_result_x[31:0]);
	always @(*) begin
		i0_predict_newp_d = dec_i0_predict_p_d;
		i0_predict_newp_d[53] = dec_i0_pc_d[1];
	end
	assign exu_pmu_i0_br_misp = i0_pp_r[55];
	assign exu_pmu_i0_br_ataken = i0_pp_r[54];
	assign exu_pmu_i0_pc4 = i0_pp_r[52];
	assign i0_valid_d = (i0_predict_p_d[37] & dec_i0_alu_decode_d) & ~dec_tlu_flush_lower_r;
	assign i0_taken_d = i0_predict_p_d[54] & dec_i0_alu_decode_d;
	generate
		if (pt[2130-:5] == 1) begin
			assign ghr_d_ns[pt[2236-:8] - 1:0] = (({pt[2236-:8] {~dec_tlu_flush_lower_r & i0_valid_d}} & {ghr_d[pt[2236-:8] - 2:0], i0_taken_d}) | ({pt[2236-:8] {~dec_tlu_flush_lower_r & ~i0_valid_d}} & ghr_d[pt[2236-:8] - 1:0])) | ({pt[2236-:8] {dec_tlu_flush_lower_r}} & ghr_x[pt[2236-:8] - 1:0]);
			assign ghr_x_ns[pt[2236-:8] - 1:0] = ({pt[2236-:8] {i0_valid_x}} & {ghr_x[pt[2236-:8] - 2:0], i0_taken_x}) | ({pt[2236-:8] {~i0_valid_x}} & ghr_x[pt[2236-:8] - 1:0]);
			assign exu_i0_br_valid_r = i0_pp_r[37];
			assign exu_i0_br_mp_r = i0_pp_r[55];
			assign exu_i0_br_way_r = i0_pp_r[32];
			assign exu_i0_br_hist_r[1:0] = {2 {i0_pp_r[37]}} & i0_pp_r[51:50];
			assign exu_i0_br_error_r = i0_pp_r[36];
			assign exu_i0_br_middle_r = i0_pp_r[52] ^ i0_pp_r[53];
			assign exu_i0_br_start_error_r = i0_pp_r[35];
			assign {exu_i0_br_fghr_r[pt[2236-:8] - 1:0], exu_i0_br_index_r[pt[2172-:9]:pt[2163-:6]]} = predpipe_r[PREDPIPESIZE - 1:pt[2139-:9]];
			assign final_predict_mp = (i0_flush_upper_x ? i0_predict_p_x : {56 {1'sb0}});
			assign final_predpipe_mp[PREDPIPESIZE - 1:0] = (i0_flush_upper_x ? predpipe_x : {PREDPIPESIZE {1'sb0}});
			assign after_flush_eghr[pt[2236-:8] - 1:0] = (i0_flush_upper_x & ~dec_tlu_flush_lower_r ? ghr_d[pt[2236-:8] - 1:0] : ghr_x[pt[2236-:8] - 1:0]);
			assign exu_mp_pkt[37] = final_predict_mp[37];
			assign exu_mp_pkt[32] = final_predict_mp[32];
			assign exu_mp_pkt[55] = final_predict_mp[55];
			assign exu_mp_pkt[34] = final_predict_mp[34];
			assign exu_mp_pkt[33] = final_predict_mp[33];
			assign exu_mp_pkt[31] = final_predict_mp[31];
			assign exu_mp_pkt[54] = final_predict_mp[54];
			assign exu_mp_pkt[53] = final_predict_mp[53];
			assign exu_mp_pkt[52] = final_predict_mp[52];
			assign exu_mp_pkt[51:50] = final_predict_mp[51:50];
			assign exu_mp_pkt[49:38] = final_predict_mp[49:38];
			assign exu_mp_fghr[pt[2236-:8] - 1:0] = after_flush_eghr[pt[2236-:8] - 1:0];
			assign {exu_mp_index[pt[2172-:9]:pt[2163-:6]], exu_mp_btag[pt[2139-:9] - 1:0]} = final_predpipe_mp[(PREDPIPESIZE - pt[2236-:8]) - 1:0];
			assign exu_mp_eghr[pt[2236-:8] - 1:0] = final_predpipe_mp[PREDPIPESIZE - 1:((pt[2172-:9] - pt[2163-:6]) + pt[2139-:9]) + 1];
		end
		else begin
			assign ghr_d_ns = {pt[2236-:8] {1'sb0}};
			assign ghr_x_ns = {pt[2236-:8] {1'sb0}};
			assign exu_mp_pkt = {56 {1'sb0}};
			assign exu_mp_eghr = {pt[2236-:8] {1'sb0}};
			assign exu_mp_fghr = {pt[2236-:8] {1'sb0}};
			assign exu_mp_index = {(pt[2172-:9] >= pt[2163-:6] ? (pt[2172-:9] - pt[2163-:6]) + 1 : (pt[2163-:6] - pt[2172-:9]) + 1) {1'sb0}};
			assign exu_mp_btag = {pt[2139-:9] {1'sb0}};
			assign exu_i0_br_hist_r = {2 {1'sb0}};
			assign exu_i0_br_error_r = 1'b0;
			assign exu_i0_br_start_error_r = 1'b0;
			assign exu_i0_br_index_r = {(pt[2172-:9] >= pt[2163-:6] ? (pt[2172-:9] - pt[2163-:6]) + 1 : (pt[2163-:6] - pt[2172-:9]) + 1) {1'sb0}};
			assign exu_i0_br_valid_r = 1'b0;
			assign exu_i0_br_mp_r = 1'b0;
			assign exu_i0_br_middle_r = 1'b0;
			assign exu_i0_br_fghr_r = {pt[2236-:8] {1'sb0}};
			assign exu_i0_br_way_r = 1'b0;
		end
	endgenerate
	assign exu_flush_path_final[31:1] = ({31 {dec_tlu_flush_lower_r}} & dec_tlu_flush_path_r[31:1]) | ({31 {~dec_tlu_flush_lower_r & i0_flush_upper_d}} & i0_flush_path_d[31:1]);
	assign exu_npc_r[31:1] = (i0_pred_correct_upper_r ? pred_correct_npc_r[31:1] : i0_flush_path_upper_r[31:1]);
endmodule
module eb1_dma_ctrl (
	clk,
	free_clk,
	rst_l,
	dma_bus_clk_en,
	clk_override,
	scan_mode,
	dbg_cmd_addr,
	dbg_cmd_wrdata,
	dbg_cmd_valid,
	dbg_cmd_write,
	dbg_cmd_type,
	dbg_cmd_size,
	dbg_dma_bubble,
	dma_dbg_ready,
	dma_dbg_cmd_done,
	dma_dbg_cmd_fail,
	dma_dbg_rddata,
	dma_dccm_req,
	dma_iccm_req,
	dma_mem_tag,
	dma_mem_addr,
	dma_mem_sz,
	dma_mem_write,
	dma_mem_wdata,
	dccm_dma_rvalid,
	dccm_dma_ecc_error,
	dccm_dma_rtag,
	dccm_dma_rdata,
	iccm_dma_rvalid,
	iccm_dma_ecc_error,
	iccm_dma_rtag,
	iccm_dma_rdata,
	dma_active,
	dma_dccm_stall_any,
	dma_iccm_stall_any,
	dccm_ready,
	iccm_ready,
	dec_tlu_dma_qos_prty,
	dma_pmu_dccm_read,
	dma_pmu_dccm_write,
	dma_pmu_any_read,
	dma_pmu_any_write,
	dma_axi_awvalid,
	dma_axi_awready,
	dma_axi_awid,
	dma_axi_awaddr,
	dma_axi_awsize,
	dma_axi_wvalid,
	dma_axi_wready,
	dma_axi_wdata,
	dma_axi_wstrb,
	dma_axi_bvalid,
	dma_axi_bready,
	dma_axi_bresp,
	dma_axi_bid,
	dma_axi_arvalid,
	dma_axi_arready,
	dma_axi_arid,
	dma_axi_araddr,
	dma_axi_arsize,
	dma_axi_rvalid,
	dma_axi_rready,
	dma_axi_rid,
	dma_axi_rdata,
	dma_axi_rresp,
	dma_axi_rlast
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire free_clk;
	input wire rst_l;
	input wire dma_bus_clk_en;
	input wire clk_override;
	input wire scan_mode;
	input wire [31:0] dbg_cmd_addr;
	input wire [31:0] dbg_cmd_wrdata;
	input wire dbg_cmd_valid;
	input wire dbg_cmd_write;
	input wire [1:0] dbg_cmd_type;
	input wire [1:0] dbg_cmd_size;
	input wire dbg_dma_bubble;
	output wire dma_dbg_ready;
	output wire dma_dbg_cmd_done;
	output wire dma_dbg_cmd_fail;
	output wire [31:0] dma_dbg_rddata;
	output wire dma_dccm_req;
	output wire dma_iccm_req;
	output wire [2:0] dma_mem_tag;
	output wire [31:0] dma_mem_addr;
	output wire [2:0] dma_mem_sz;
	output wire dma_mem_write;
	output wire [63:0] dma_mem_wdata;
	input wire dccm_dma_rvalid;
	input wire dccm_dma_ecc_error;
	input wire [2:0] dccm_dma_rtag;
	input wire [63:0] dccm_dma_rdata;
	input wire iccm_dma_rvalid;
	input wire iccm_dma_ecc_error;
	input wire [2:0] iccm_dma_rtag;
	input wire [63:0] iccm_dma_rdata;
	output wire dma_active;
	output wire dma_dccm_stall_any;
	output wire dma_iccm_stall_any;
	input wire dccm_ready;
	input wire iccm_ready;
	input wire [2:0] dec_tlu_dma_qos_prty;
	output wire dma_pmu_dccm_read;
	output wire dma_pmu_dccm_write;
	output wire dma_pmu_any_read;
	output wire dma_pmu_any_write;
	input wire dma_axi_awvalid;
	output wire dma_axi_awready;
	input wire [pt[1235-:8] - 1:0] dma_axi_awid;
	input wire [31:0] dma_axi_awaddr;
	input wire [2:0] dma_axi_awsize;
	input wire dma_axi_wvalid;
	output wire dma_axi_wready;
	input wire [63:0] dma_axi_wdata;
	input wire [7:0] dma_axi_wstrb;
	output wire dma_axi_bvalid;
	input wire dma_axi_bready;
	output wire [1:0] dma_axi_bresp;
	output wire [pt[1235-:8] - 1:0] dma_axi_bid;
	input wire dma_axi_arvalid;
	output wire dma_axi_arready;
	input wire [pt[1235-:8] - 1:0] dma_axi_arid;
	input wire [31:0] dma_axi_araddr;
	input wire [2:0] dma_axi_arsize;
	output wire dma_axi_rvalid;
	input wire dma_axi_rready;
	output wire [pt[1235-:8] - 1:0] dma_axi_rid;
	output wire [63:0] dma_axi_rdata;
	output wire [1:0] dma_axi_rresp;
	output wire dma_axi_rlast;
	localparam DEPTH = pt[1257-:7];
	localparam DEPTH_PTR = $clog2(DEPTH);
	localparam NACK_COUNT = 7;
	wire [DEPTH - 1:0] fifo_valid;
	wire [(DEPTH * 2) - 1:0] fifo_error;
	wire [DEPTH - 1:0] fifo_error_bus;
	wire [DEPTH - 1:0] fifo_rpend;
	wire [DEPTH - 1:0] fifo_done;
	wire [DEPTH - 1:0] fifo_done_bus;
	wire [(DEPTH * 32) - 1:0] fifo_addr;
	wire [(DEPTH * 3) - 1:0] fifo_sz;
	wire [(DEPTH * 8) - 1:0] fifo_byteen;
	wire [DEPTH - 1:0] fifo_write;
	wire [DEPTH - 1:0] fifo_posted_write;
	wire [DEPTH - 1:0] fifo_dbg;
	wire [(DEPTH * 64) - 1:0] fifo_data;
	wire [(DEPTH * pt[1235-:8]) - 1:0] fifo_tag;
	wire [(DEPTH * pt[1250-:9]) - 1:0] fifo_mid;
	wire [(DEPTH * pt[1241-:6]) - 1:0] fifo_prty;
	wire [DEPTH - 1:0] fifo_cmd_en;
	wire [DEPTH - 1:0] fifo_data_en;
	wire [DEPTH - 1:0] fifo_pend_en;
	wire [DEPTH - 1:0] fifo_done_en;
	wire [DEPTH - 1:0] fifo_done_bus_en;
	wire [DEPTH - 1:0] fifo_error_en;
	wire [DEPTH - 1:0] fifo_error_bus_en;
	wire [DEPTH - 1:0] fifo_reset;
	wire [(DEPTH * 2) - 1:0] fifo_error_in;
	wire [(DEPTH * 64) - 1:0] fifo_data_in;
	wire fifo_write_in;
	wire fifo_posted_write_in;
	wire fifo_dbg_in;
	wire [31:0] fifo_addr_in;
	wire [2:0] fifo_sz_in;
	wire [7:0] fifo_byteen_in;
	wire [DEPTH_PTR - 1:0] RspPtr;
	wire [DEPTH_PTR - 1:0] NxtRspPtr;
	wire [DEPTH_PTR - 1:0] WrPtr;
	wire [DEPTH_PTR - 1:0] NxtWrPtr;
	wire [DEPTH_PTR - 1:0] RdPtr;
	wire [DEPTH_PTR - 1:0] NxtRdPtr;
	wire WrPtrEn;
	wire RdPtrEn;
	wire RspPtrEn;
	wire [1:0] dma_dbg_sz;
	wire [1:0] dma_dbg_addr;
	wire [31:0] dma_dbg_mem_rddata;
	wire [31:0] dma_dbg_mem_wrdata;
	wire dma_dbg_cmd_error;
	wire dma_dbg_cmd_done_q;
	wire fifo_full;
	wire fifo_full_spec;
	wire fifo_empty;
	wire dma_address_error;
	wire dma_alignment_error;
	reg [3:0] num_fifo_vld;
	wire dma_mem_req;
	wire [31:0] dma_mem_addr_int;
	wire [2:0] dma_mem_sz_int;
	wire [7:0] dma_mem_byteen;
	wire dma_mem_addr_in_dccm;
	wire dma_mem_addr_in_iccm;
	wire dma_mem_addr_in_pic;
	wire dma_mem_addr_in_pic_region_nc;
	wire dma_mem_addr_in_dccm_region_nc;
	wire dma_mem_addr_in_iccm_region_nc;
	wire [2:0] dma_nack_count;
	wire [2:0] dma_nack_count_d;
	wire [2:0] dma_nack_count_csr;
	wire dma_buffer_c1_clken;
	wire dma_free_clken;
	wire dma_buffer_c1_clk;
	wire dma_free_clk;
	wire dma_bus_clk;
	wire bus_rsp_valid;
	wire bus_rsp_sent;
	wire bus_cmd_valid;
	wire bus_cmd_sent;
	wire bus_cmd_write;
	wire bus_cmd_posted_write;
	wire [7:0] bus_cmd_byteen;
	wire [2:0] bus_cmd_sz;
	wire [31:0] bus_cmd_addr;
	wire [63:0] bus_cmd_wdata;
	wire [pt[1235-:8] - 1:0] bus_cmd_tag;
	wire [pt[1250-:9] - 1:0] bus_cmd_mid;
	wire [pt[1241-:6] - 1:0] bus_cmd_prty;
	wire bus_posted_write_done;
	wire fifo_full_spec_bus;
	wire dbg_dma_bubble_bus;
	wire stall_dma_in;
	wire dma_fifo_ready;
	wire wrbuf_en;
	wire wrbuf_data_en;
	wire wrbuf_cmd_sent;
	wire wrbuf_rst;
	wire wrbuf_data_rst;
	wire wrbuf_vld;
	wire wrbuf_data_vld;
	wire [pt[1235-:8] - 1:0] wrbuf_tag;
	wire [2:0] wrbuf_sz;
	wire [31:0] wrbuf_addr;
	wire [63:0] wrbuf_data;
	wire [7:0] wrbuf_byteen;
	wire rdbuf_en;
	wire rdbuf_cmd_sent;
	wire rdbuf_rst;
	wire rdbuf_vld;
	wire [pt[1235-:8] - 1:0] rdbuf_tag;
	wire [2:0] rdbuf_sz;
	wire [31:0] rdbuf_addr;
	wire axi_mstr_prty_in;
	wire axi_mstr_prty_en;
	wire axi_mstr_priority;
	wire axi_mstr_sel;
	wire axi_rsp_valid;
	wire axi_rsp_sent;
	wire axi_rsp_write;
	wire [pt[1235-:8] - 1:0] axi_rsp_tag;
	wire [1:0] axi_rsp_error;
	wire [63:0] axi_rsp_rdata;
	assign fifo_addr_in[31:0] = (dbg_cmd_valid ? dbg_cmd_addr[31:0] : bus_cmd_addr[31:0]);
	assign fifo_byteen_in[7:0] = {8 {~dbg_cmd_valid}} & bus_cmd_byteen[7:0];
	assign fifo_sz_in[2:0] = (dbg_cmd_valid ? {1'b0, dbg_cmd_size[1:0]} : bus_cmd_sz[2:0]);
	assign fifo_write_in = (dbg_cmd_valid ? dbg_cmd_write : bus_cmd_write);
	assign fifo_posted_write_in = ~dbg_cmd_valid & bus_cmd_posted_write;
	assign fifo_dbg_in = dbg_cmd_valid;
	generate
		genvar i;
		for (i = 0; i < DEPTH; i = i + 1) begin : GenFifo
			assign fifo_cmd_en[i] = ((bus_cmd_sent & dma_bus_clk_en) | (dbg_cmd_valid & dbg_cmd_type[1])) & (i == WrPtr[DEPTH_PTR - 1:0]);
			function automatic [DEPTH_PTR - 1:0] sv2v_cast_87E0F;
				input reg [DEPTH_PTR - 1:0] inp;
				sv2v_cast_87E0F = inp;
			endfunction
			assign fifo_data_en[i] = ((((((bus_cmd_sent & fifo_write_in) & dma_bus_clk_en) | ((dbg_cmd_valid & dbg_cmd_type[1]) & dbg_cmd_write)) & (i == WrPtr[DEPTH_PTR - 1:0])) | ((dma_address_error | dma_alignment_error) & (i == RdPtr[DEPTH_PTR - 1:0]))) | (dccm_dma_rvalid & (i == sv2v_cast_87E0F(dccm_dma_rtag[2:0])))) | (iccm_dma_rvalid & (i == sv2v_cast_87E0F(iccm_dma_rtag[2:0])));
			assign fifo_pend_en[i] = ((dma_dccm_req | dma_iccm_req) & ~dma_mem_write) & (i == RdPtr[DEPTH_PTR - 1:0]);
			assign fifo_error_en[i] = ((((dma_address_error | dma_alignment_error) | dma_dbg_cmd_error) & (i == RdPtr[DEPTH_PTR - 1:0])) | ((dccm_dma_rvalid & dccm_dma_ecc_error) & (i == sv2v_cast_87E0F(dccm_dma_rtag[2:0])))) | ((iccm_dma_rvalid & iccm_dma_ecc_error) & (i == sv2v_cast_87E0F(iccm_dma_rtag[2:0])));
			assign fifo_error_bus_en[i] = ((|fifo_error_in[(i * 2) + 1-:2] & fifo_error_en[i]) | |fifo_error[i * 2+:2]) & dma_bus_clk_en;
			assign fifo_done_en[i] = ((((|fifo_error[i * 2+:2] | fifo_error_en[i]) | ((dma_dccm_req | dma_iccm_req) & dma_mem_write)) & (i == RdPtr[DEPTH_PTR - 1:0])) | (dccm_dma_rvalid & (i == sv2v_cast_87E0F(dccm_dma_rtag[2:0])))) | (iccm_dma_rvalid & (i == sv2v_cast_87E0F(iccm_dma_rtag[2:0])));
			assign fifo_done_bus_en[i] = (fifo_done_en[i] | fifo_done[i]) & dma_bus_clk_en;
			assign fifo_reset[i] = (((bus_rsp_sent | bus_posted_write_done) & dma_bus_clk_en) | dma_dbg_cmd_done) & (i == RspPtr[DEPTH_PTR - 1:0]);
			assign fifo_error_in[i * 2+:2] = (dccm_dma_rvalid & (i == sv2v_cast_87E0F(dccm_dma_rtag[2:0])) ? {1'b0, dccm_dma_ecc_error} : (iccm_dma_rvalid & (i == sv2v_cast_87E0F(iccm_dma_rtag[2:0])) ? {1'b0, iccm_dma_ecc_error} : {(dma_address_error | dma_alignment_error) | dma_dbg_cmd_error, dma_alignment_error}));
			assign fifo_data_in[i * 64+:64] = (fifo_error_en[i] & |fifo_error_in[i * 2+:2] ? {32'b00000000000000000000000000000000, fifo_addr[i * 32+:32]} : (dccm_dma_rvalid & (i == sv2v_cast_87E0F(dccm_dma_rtag[2:0])) ? dccm_dma_rdata[63:0] : (iccm_dma_rvalid & (i == sv2v_cast_87E0F(iccm_dma_rtag[2:0])) ? iccm_dma_rdata[63:0] : (dbg_cmd_valid ? {2 {dma_dbg_mem_wrdata[31:0]}} : bus_cmd_wdata[63:0]))));
			rvdffsc #(.WIDTH(1)) fifo_valid_dff(
				.din(1'b1),
				.dout(fifo_valid[i]),
				.en(fifo_cmd_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffsc #(.WIDTH(2)) fifo_error_dff(
				.din(fifo_error_in[i * 2+:2]),
				.dout(fifo_error[i * 2+:2]),
				.en(fifo_error_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffsc #(.WIDTH(1)) fifo_error_bus_dff(
				.din(1'b1),
				.dout(fifo_error_bus[i]),
				.en(fifo_error_bus_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffsc #(.WIDTH(1)) fifo_rpend_dff(
				.din(1'b1),
				.dout(fifo_rpend[i]),
				.en(fifo_pend_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffsc #(.WIDTH(1)) fifo_done_dff(
				.din(1'b1),
				.dout(fifo_done[i]),
				.en(fifo_done_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffsc #(.WIDTH(1)) fifo_done_bus_dff(
				.din(1'b1),
				.dout(fifo_done_bus[i]),
				.en(fifo_done_bus_en[i]),
				.clear(fifo_reset[i]),
				.clk(dma_free_clk),
				.rst_l(rst_l)
			);
			rvdffe #(.WIDTH(32)) fifo_addr_dff(
				.din(fifo_addr_in[31:0]),
				.dout(fifo_addr[i * 32+:32]),
				.en(fifo_cmd_en[i]),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
			rvdffs #(.WIDTH(3)) fifo_sz_dff(
				.din(fifo_sz_in[2:0]),
				.dout(fifo_sz[i * 3+:3]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(8)) fifo_byteen_dff(
				.din(fifo_byteen_in[7:0]),
				.dout(fifo_byteen[i * 8+:8]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) fifo_write_dff(
				.din(fifo_write_in),
				.dout(fifo_write[i]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) fifo_posted_write_dff(
				.din(fifo_posted_write_in),
				.dout(fifo_posted_write[i]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) fifo_dbg_dff(
				.din(fifo_dbg_in),
				.dout(fifo_dbg[i]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffe #(.WIDTH(64)) fifo_data_dff(
				.din(fifo_data_in[i * 64+:64]),
				.dout(fifo_data[i * 64+:64]),
				.en(fifo_data_en[i]),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
			rvdffs #(.WIDTH(pt[1235-:8])) fifo_tag_dff(
				.din(bus_cmd_tag[pt[1235-:8] - 1:0]),
				.dout(fifo_tag[(i * pt[1235-:8]) + (pt[1235-:8] - 1)-:pt[1235-:8]]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(pt[1250-:9])) fifo_mid_dff(
				.din(bus_cmd_mid[pt[1250-:9] - 1:0]),
				.dout(fifo_mid[(i * pt[1250-:9]) + (pt[1250-:9] - 1)-:pt[1250-:9]]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(pt[1241-:6])) fifo_prty_dff(
				.din(bus_cmd_prty[pt[1241-:6] - 1:0]),
				.dout(fifo_prty[(i * pt[1241-:6]) + (pt[1241-:6] - 1)-:pt[1241-:6]]),
				.en(fifo_cmd_en[i]),
				.clk(dma_buffer_c1_clk),
				.rst_l(rst_l)
			);
		end
	endgenerate
	assign NxtWrPtr[DEPTH_PTR - 1:0] = (WrPtr[DEPTH_PTR - 1:0] == (DEPTH - 1) ? {DEPTH_PTR {1'sb0}} : WrPtr[DEPTH_PTR - 1:0] + 1'b1);
	assign NxtRdPtr[DEPTH_PTR - 1:0] = (RdPtr[DEPTH_PTR - 1:0] == (DEPTH - 1) ? {DEPTH_PTR {1'sb0}} : RdPtr[DEPTH_PTR - 1:0] + 1'b1);
	assign NxtRspPtr[DEPTH_PTR - 1:0] = (RspPtr[DEPTH_PTR - 1:0] == (DEPTH - 1) ? {DEPTH_PTR {1'sb0}} : RspPtr[DEPTH_PTR - 1:0] + 1'b1);
	assign WrPtrEn = |fifo_cmd_en[DEPTH - 1:0];
	assign RdPtrEn = (dma_dccm_req | dma_iccm_req) | ((dma_address_error | dma_alignment_error) | dma_dbg_cmd_error);
	assign RspPtrEn = dma_dbg_cmd_done | ((bus_rsp_sent | bus_posted_write_done) & dma_bus_clk_en);
	rvdffs #(.WIDTH(DEPTH_PTR)) WrPtr_dff(
		.din(NxtWrPtr[DEPTH_PTR - 1:0]),
		.dout(WrPtr[DEPTH_PTR - 1:0]),
		.en(WrPtrEn),
		.clk(dma_free_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(DEPTH_PTR)) RdPtr_dff(
		.din(NxtRdPtr[DEPTH_PTR - 1:0]),
		.dout(RdPtr[DEPTH_PTR - 1:0]),
		.en(RdPtrEn),
		.clk(dma_free_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(DEPTH_PTR)) RspPtr_dff(
		.din(NxtRspPtr[DEPTH_PTR - 1:0]),
		.dout(RspPtr[DEPTH_PTR - 1:0]),
		.en(RspPtrEn),
		.clk(dma_free_clk),
		.rst_l(rst_l)
	);
	assign fifo_full = fifo_full_spec_bus;
	always @(*) begin
		num_fifo_vld[3:0] = {3'b000, bus_cmd_sent} - {3'b000, bus_rsp_sent};
		begin : sv2v_autoblock_41
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				num_fifo_vld[3:0] = num_fifo_vld[3:0] + {3'b000, fifo_valid[i]};
		end
	end
	assign fifo_full_spec = num_fifo_vld[3:0] >= DEPTH;
	assign dma_fifo_ready = ~(fifo_full | dbg_dma_bubble_bus);
	assign dma_address_error = ((fifo_valid[RdPtr] & ~fifo_done[RdPtr]) & ~fifo_dbg[RdPtr]) & ~(dma_mem_addr_in_dccm | dma_mem_addr_in_iccm);
	assign dma_alignment_error = (((fifo_valid[RdPtr] & ~fifo_done[RdPtr]) & ~fifo_dbg[RdPtr]) & ~dma_address_error) & ((((((((dma_mem_sz_int[2:0] == 3'h1) & dma_mem_addr_int[0]) | ((dma_mem_sz_int[2:0] == 3'h2) & |dma_mem_addr_int[1:0])) | ((dma_mem_sz_int[2:0] == 3'h3) & |dma_mem_addr_int[2:0])) | (dma_mem_addr_in_iccm & ~((dma_mem_sz_int[1:0] == 2'b10) | (dma_mem_sz_int[1:0] == 2'b11)))) | ((dma_mem_addr_in_dccm & dma_mem_write) & ~((dma_mem_sz_int[1:0] == 2'b10) | (dma_mem_sz_int[1:0] == 2'b11)))) | ((dma_mem_write & (dma_mem_sz_int[2:0] == 3'h2)) & (dma_mem_byteen[dma_mem_addr_int[2:0]+:4] != 4'hf))) | ((dma_mem_write & (dma_mem_sz_int[2:0] == 3'h3)) & ~(((dma_mem_byteen[7:0] == 8'h0f) | (dma_mem_byteen[7:0] == 8'hf0)) | (dma_mem_byteen[7:0] == 8'hff))));
	assign dma_dbg_ready = fifo_empty & dbg_dma_bubble;
	assign dma_dbg_cmd_done = (fifo_valid[RspPtr] & fifo_dbg[RspPtr]) & fifo_done[RspPtr];
	assign dma_dbg_cmd_fail = |fifo_error[RspPtr * 2+:2];
	assign dma_dbg_sz[1:0] = fifo_sz[(RspPtr * 3) + 1-:2];
	assign dma_dbg_addr[1:0] = fifo_addr[(RspPtr * 32) + 1-:2];
	assign dma_dbg_mem_rddata[31:0] = (fifo_addr[(RspPtr * 32) + 2] ? fifo_data[(RspPtr * 64) + 63-:32] : fifo_data[(RspPtr * 64) + 31-:32]);
	assign dma_dbg_rddata[31:0] = (({32 {dma_dbg_sz[1:0] == 2'h0}} & ((dma_dbg_mem_rddata[31:0] >> (8 * dma_dbg_addr[1:0])) & 32'h000000ff)) | ({32 {dma_dbg_sz[1:0] == 2'h1}} & ((dma_dbg_mem_rddata[31:0] >> (16 * dma_dbg_addr[1])) & 32'h0000ffff))) | ({32 {dma_dbg_sz[1:0] == 2'h2}} & dma_dbg_mem_rddata[31:0]);
	assign dma_dbg_cmd_error = ((fifo_valid[RdPtr] & ~fifo_done[RdPtr]) & fifo_dbg[RdPtr]) & (~((dma_mem_addr_in_dccm | dma_mem_addr_in_iccm) | dma_mem_addr_in_pic) | ((dma_mem_addr_in_iccm | dma_mem_addr_in_pic) & (dma_mem_sz_int[1:0] != 2'b10)));
	assign dma_dbg_mem_wrdata[31:0] = (({32 {dbg_cmd_size[1:0] == 2'h0}} & {4 {dbg_cmd_wrdata[7:0]}}) | ({32 {dbg_cmd_size[1:0] == 2'h1}} & {2 {dbg_cmd_wrdata[15:0]}})) | ({32 {dbg_cmd_size[1:0] == 2'h2}} & dbg_cmd_wrdata[31:0]);
	assign dma_dccm_stall_any = (dma_mem_req & (dma_mem_addr_in_dccm | dma_mem_addr_in_pic)) & (dma_nack_count >= dma_nack_count_csr);
	assign dma_iccm_stall_any = (dma_mem_req & dma_mem_addr_in_iccm) & (dma_nack_count >= dma_nack_count_csr);
	assign fifo_empty = ~(|fifo_valid[DEPTH - 1:0] | bus_cmd_sent);
	assign dma_nack_count_csr[2:0] = dec_tlu_dma_qos_prty[2:0];
	assign dma_nack_count_d[2:0] = (dma_nack_count[2:0] >= dma_nack_count_csr[2:0] ? {3 {~(dma_dccm_req | dma_iccm_req)}} & dma_nack_count[2:0] : (dma_mem_req & ~(dma_dccm_req | dma_iccm_req) ? dma_nack_count[2:0] + 1'b1 : 3'b000));
	rvdffs #(.WIDTH(3)) nack_count_dff(
		.din(dma_nack_count_d[2:0]),
		.dout(dma_nack_count[2:0]),
		.en(dma_mem_req),
		.clk(dma_free_clk),
		.rst_l(rst_l)
	);
	assign dma_mem_req = ((fifo_valid[RdPtr] & ~fifo_rpend[RdPtr]) & ~fifo_done[RdPtr]) & ~((dma_address_error | dma_alignment_error) | dma_dbg_cmd_error);
	assign dma_dccm_req = (dma_mem_req & (dma_mem_addr_in_dccm | dma_mem_addr_in_pic)) & dccm_ready;
	assign dma_iccm_req = (dma_mem_req & dma_mem_addr_in_iccm) & iccm_ready;
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	assign dma_mem_tag[2:0] = sv2v_cast_3(RdPtr);
	assign dma_mem_addr_int[31:0] = fifo_addr[RdPtr * 32+:32];
	assign dma_mem_sz_int[2:0] = fifo_sz[RdPtr * 3+:3];
	assign dma_mem_addr[31:0] = ((dma_mem_write & ~fifo_dbg[RdPtr]) & (dma_mem_byteen[7:0] == 8'hf0) ? {dma_mem_addr_int[31:3], 1'b1, dma_mem_addr_int[1:0]} : dma_mem_addr_int[31:0]);
	assign dma_mem_sz[2:0] = ((dma_mem_write & ~fifo_dbg[RdPtr]) & ((dma_mem_byteen[7:0] == 8'h0f) | (dma_mem_byteen[7:0] == 8'hf0)) ? 3'h2 : dma_mem_sz_int[2:0]);
	assign dma_mem_byteen[7:0] = fifo_byteen[RdPtr * 8+:8];
	assign dma_mem_write = fifo_write[RdPtr];
	assign dma_mem_wdata[63:0] = fifo_data[RdPtr * 64+:64];
	assign dma_pmu_dccm_read = dma_dccm_req & ~dma_mem_write;
	assign dma_pmu_dccm_write = dma_dccm_req & dma_mem_write;
	assign dma_pmu_any_read = (dma_dccm_req | dma_iccm_req) & ~dma_mem_write;
	assign dma_pmu_any_write = (dma_dccm_req | dma_iccm_req) & dma_mem_write;
	generate
		if (pt[1365-:5]) begin : Gen_dccm_enable
			rvrangecheck #(
				.CCM_SADR(pt[1325-:36]),
				.CCM_SIZE(pt[1289-:14])
			) addr_dccm_rangecheck(
				.addr(dma_mem_addr_int[31:0]),
				.in_range(dma_mem_addr_in_dccm),
				.in_region(dma_mem_addr_in_dccm_region_nc)
			);
		end
		else begin : Gen_dccm_disable
			assign dma_mem_addr_in_dccm = 1'b0;
			assign dma_mem_addr_in_dccm_region_nc = 1'b0;
		end
	endgenerate
	generate
		if (pt[927-:5]) begin : Gen_iccm_enable
			rvrangecheck #(
				.CCM_SADR(pt[887-:36]),
				.CCM_SIZE(pt[851-:14])
			) addr_iccm_rangecheck(
				.addr(dma_mem_addr_int[31:0]),
				.in_range(dma_mem_addr_in_iccm),
				.in_region(dma_mem_addr_in_iccm_region_nc)
			);
		end
		else begin : Gen_iccm_disable
			assign dma_mem_addr_in_iccm = 1'b0;
			assign dma_mem_addr_in_iccm_region_nc = 1'b0;
		end
	endgenerate
	rvrangecheck #(
		.CCM_SADR(pt[130-:36]),
		.CCM_SIZE(pt[69-:13])
	) addr_pic_rangecheck(
		.addr(dma_mem_addr_int[31:0]),
		.in_range(dma_mem_addr_in_pic),
		.in_region(dma_mem_addr_in_pic_region_nc)
	);
	rvdff_fpga #(.WIDTH(1)) fifo_full_bus_ff(
		.din(fifo_full_spec),
		.dout(fifo_full_spec_bus),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) dbg_dma_bubble_ff(
		.din(dbg_dma_bubble),
		.dout(dbg_dma_bubble_bus),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) dma_dbg_cmd_doneff(
		.din(dma_dbg_cmd_done),
		.dout(dma_dbg_cmd_done_q),
		.clk(free_clk),
		.rst_l(rst_l)
	);
	assign dma_buffer_c1_clken = ((bus_cmd_valid & dma_bus_clk_en) | dbg_cmd_valid) | clk_override;
	assign dma_free_clken = (((((bus_cmd_valid | bus_rsp_valid) | dbg_cmd_valid) | dma_dbg_cmd_done) | dma_dbg_cmd_done_q) | |fifo_valid[DEPTH - 1:0]) | clk_override;
	rvoclkhdr dma_buffer_c1cgc(
		.en(dma_buffer_c1_clken),
		.l1clk(dma_buffer_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr dma_free_cgc(
		.en(dma_free_clken),
		.l1clk(dma_free_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr dma_bus_cgc(
		.en(dma_bus_clk_en),
		.l1clk(dma_bus_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign wrbuf_en = dma_axi_awvalid & dma_axi_awready;
	assign wrbuf_data_en = dma_axi_wvalid & dma_axi_wready;
	assign wrbuf_cmd_sent = bus_cmd_sent & bus_cmd_write;
	assign wrbuf_rst = wrbuf_cmd_sent & ~wrbuf_en;
	assign wrbuf_data_rst = wrbuf_cmd_sent & ~wrbuf_data_en;
	rvdffsc_fpga #(.WIDTH(1)) wrbuf_vldff(
		.din(1'b1),
		.dout(wrbuf_vld),
		.en(wrbuf_en),
		.clear(wrbuf_rst),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffsc_fpga #(.WIDTH(1)) wrbuf_data_vldff(
		.din(1'b1),
		.dout(wrbuf_data_vld),
		.en(wrbuf_data_en),
		.clear(wrbuf_data_rst),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(pt[1235-:8])) wrbuf_tagff(
		.din(dma_axi_awid[pt[1235-:8] - 1:0]),
		.dout(wrbuf_tag[pt[1235-:8] - 1:0]),
		.en(wrbuf_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(3)) wrbuf_szff(
		.din(dma_axi_awsize[2:0]),
		.dout(wrbuf_sz[2:0]),
		.en(wrbuf_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) wrbuf_addrff(
		.din(dma_axi_awaddr[31:0]),
		.dout(wrbuf_addr[31:0]),
		.en(wrbuf_en & dma_bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffe #(.WIDTH(64)) wrbuf_dataff(
		.din(dma_axi_wdata[63:0]),
		.dout(wrbuf_data[63:0]),
		.en(wrbuf_data_en & dma_bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffs_fpga #(.WIDTH(8)) wrbuf_byteenff(
		.din(dma_axi_wstrb[7:0]),
		.dout(wrbuf_byteen[7:0]),
		.en(wrbuf_data_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	assign rdbuf_en = dma_axi_arvalid & dma_axi_arready;
	assign rdbuf_cmd_sent = bus_cmd_sent & ~bus_cmd_write;
	assign rdbuf_rst = rdbuf_cmd_sent & ~rdbuf_en;
	rvdffsc_fpga #(.WIDTH(1)) rdbuf_vldff(
		.din(1'b1),
		.dout(rdbuf_vld),
		.en(rdbuf_en),
		.clear(rdbuf_rst),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(pt[1235-:8])) rdbuf_tagff(
		.din(dma_axi_arid[pt[1235-:8] - 1:0]),
		.dout(rdbuf_tag[pt[1235-:8] - 1:0]),
		.en(rdbuf_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(3)) rdbuf_szff(
		.din(dma_axi_arsize[2:0]),
		.dout(rdbuf_sz[2:0]),
		.en(rdbuf_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) rdbuf_addrff(
		.din(dma_axi_araddr[31:0]),
		.dout(rdbuf_addr[31:0]),
		.en(rdbuf_en & dma_bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	assign dma_axi_awready = ~(wrbuf_vld & ~wrbuf_cmd_sent);
	assign dma_axi_wready = ~(wrbuf_data_vld & ~wrbuf_cmd_sent);
	assign dma_axi_arready = ~(rdbuf_vld & ~rdbuf_cmd_sent);
	assign bus_cmd_valid = (wrbuf_vld & wrbuf_data_vld) | rdbuf_vld;
	assign bus_cmd_sent = bus_cmd_valid & dma_fifo_ready;
	assign bus_cmd_write = axi_mstr_sel;
	assign bus_cmd_posted_write = 1'b0;
	assign bus_cmd_addr[31:0] = (axi_mstr_sel ? wrbuf_addr[31:0] : rdbuf_addr[31:0]);
	assign bus_cmd_sz[2:0] = (axi_mstr_sel ? wrbuf_sz[2:0] : rdbuf_sz[2:0]);
	assign bus_cmd_wdata[63:0] = wrbuf_data[63:0];
	assign bus_cmd_byteen[7:0] = wrbuf_byteen[7:0];
	assign bus_cmd_tag[pt[1235-:8] - 1:0] = (axi_mstr_sel ? wrbuf_tag[pt[1235-:8] - 1:0] : rdbuf_tag[pt[1235-:8] - 1:0]);
	assign bus_cmd_mid[pt[1250-:9] - 1:0] = {pt[1250-:9] {1'sb0}};
	assign bus_cmd_prty[pt[1241-:6] - 1:0] = {pt[1241-:6] {1'sb0}};
	assign axi_mstr_sel = ((wrbuf_vld & wrbuf_data_vld) & rdbuf_vld ? axi_mstr_priority : wrbuf_vld & wrbuf_data_vld);
	assign axi_mstr_prty_in = ~axi_mstr_priority;
	assign axi_mstr_prty_en = bus_cmd_sent;
	rvdffs_fpga #(.WIDTH(1)) mstr_prtyff(
		.din(axi_mstr_prty_in),
		.dout(axi_mstr_priority),
		.en(axi_mstr_prty_en),
		.clk(dma_bus_clk),
		.clken(dma_bus_clk_en),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	assign axi_rsp_valid = (fifo_valid[RspPtr] & ~fifo_dbg[RspPtr]) & fifo_done_bus[RspPtr];
	assign axi_rsp_rdata[63:0] = fifo_data[RspPtr * 64+:64];
	assign axi_rsp_write = fifo_write[RspPtr];
	assign axi_rsp_error[1:0] = (fifo_error[RspPtr * 2] ? 2'b10 : (fifo_error[(RspPtr * 2) + 1] ? 2'b11 : 2'b00));
	assign axi_rsp_tag[pt[1235-:8] - 1:0] = fifo_tag[RspPtr * pt[1235-:8]+:pt[1235-:8]];
	assign dma_axi_bvalid = axi_rsp_valid & axi_rsp_write;
	assign dma_axi_bresp[1:0] = axi_rsp_error[1:0];
	assign dma_axi_bid[pt[1235-:8] - 1:0] = axi_rsp_tag[pt[1235-:8] - 1:0];
	assign dma_axi_rvalid = axi_rsp_valid & ~axi_rsp_write;
	assign dma_axi_rresp[1:0] = axi_rsp_error;
	assign dma_axi_rdata[63:0] = axi_rsp_rdata[63:0];
	assign dma_axi_rlast = 1'b1;
	assign dma_axi_rid[pt[1235-:8] - 1:0] = axi_rsp_tag[pt[1235-:8] - 1:0];
	assign bus_posted_write_done = 1'b0;
	assign bus_rsp_valid = dma_axi_bvalid | dma_axi_rvalid;
	assign bus_rsp_sent = (dma_axi_bvalid & dma_axi_bready) | (dma_axi_rvalid & dma_axi_rready);
	assign dma_active = (wrbuf_vld | rdbuf_vld) | |fifo_valid[DEPTH - 1:0];
endmodule
module eb1_exu_alu_ctl (
	clk,
	rst_l,
	scan_mode,
	flush_upper_x,
	flush_lower_r,
	enable,
	valid_in,
	ap,
	csr_ren_in,
	csr_rddata_in,
	a_in,
	b_in,
	pc_in,
	pp_in,
	brimm_in,
	result_ff,
	flush_upper_out,
	flush_final_out,
	flush_path_out,
	pc_ff,
	pred_correct_out,
	predict_p_out
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire flush_upper_x;
	input wire flush_lower_r;
	input wire enable;
	input wire valid_in;
	input wire [43:0] ap;
	input wire csr_ren_in;
	input wire [31:0] csr_rddata_in;
	input wire signed [31:0] a_in;
	input wire [31:0] b_in;
	input wire [31:1] pc_in;
	input wire [55:0] pp_in;
	input wire [12:1] brimm_in;
	output wire [31:0] result_ff;
	output wire flush_upper_out;
	output wire flush_final_out;
	output wire [31:1] flush_path_out;
	output wire [31:1] pc_ff;
	output wire pred_correct_out;
	output reg [55:0] predict_p_out;
	wire [31:0] zba_a_in;
	wire [31:0] aout;
	wire cout;
	wire ov;
	wire neg;
	wire [31:0] lout;
	wire [31:0] sout;
	wire sel_shift;
	wire sel_adder;
	wire slt_one;
	wire actual_taken;
	wire [31:1] pcout;
	wire cond_mispredict;
	wire target_mispredict;
	wire eq;
	wire ne;
	wire lt;
	wire ge;
	wire any_jal;
	wire [1:0] newhist;
	wire sel_pc;
	wire [31:0] csr_write_data;
	wire [31:0] result;
	wire ap_clz;
	wire ap_ctz;
	wire ap_pcnt;
	wire ap_sext_b;
	wire ap_sext_h;
	wire ap_min;
	wire ap_max;
	wire ap_pack;
	wire ap_packu;
	wire ap_packh;
	wire ap_rol;
	wire ap_ror;
	wire ap_rev;
	wire ap_rev8;
	wire ap_orc_b;
	wire ap_orc16;
	wire ap_zbb;
	wire ap_sbset;
	wire ap_sbclr;
	wire ap_sbinv;
	wire ap_sbext;
	wire ap_slo;
	wire ap_sro;
	wire ap_sh1add;
	wire ap_sh2add;
	wire ap_sh3add;
	wire ap_zba;
	generate
		if (pt[2207-:5] == 1) begin
			assign ap_clz = ap[43];
			assign ap_ctz = ap[42];
			assign ap_pcnt = ap[41];
			assign ap_sext_b = ap[40];
			assign ap_sext_h = ap[39];
			assign ap_min = ap[36];
			assign ap_max = ap[35];
		end
		else begin
			assign ap_clz = 1'b0;
			assign ap_ctz = 1'b0;
			assign ap_pcnt = 1'b0;
			assign ap_sext_b = 1'b0;
			assign ap_sext_h = 1'b0;
			assign ap_min = 1'b0;
			assign ap_max = 1'b0;
		end
	endgenerate
	generate
		if ((pt[2207-:5] == 1) | (pt[2187-:5] == 1)) begin
			assign ap_pack = ap[34];
			assign ap_packu = ap[33];
			assign ap_packh = ap[32];
			assign ap_rol = ap[31];
			assign ap_ror = ap[30];
			assign ap_rev = ap[29] & (b_in[4:0] == 5'b11111);
			assign ap_rev8 = ap[29] & (b_in[4:0] == 5'b11000);
			assign ap_orc_b = ap[28] & (b_in[4:0] == 5'b00111);
			assign ap_orc16 = ap[28] & (b_in[4:0] == 5'b10000);
			assign ap_zbb = ap[27];
		end
		else begin
			assign ap_pack = 1'b0;
			assign ap_packu = 1'b0;
			assign ap_packh = 1'b0;
			assign ap_rol = 1'b0;
			assign ap_ror = 1'b0;
			assign ap_rev = 1'b0;
			assign ap_rev8 = 1'b0;
			assign ap_orc_b = 1'b0;
			assign ap_orc16 = 1'b0;
			assign ap_zbb = 1'b0;
		end
	endgenerate
	generate
		if (pt[2177-:5] == 1) begin
			assign ap_sbset = ap[26];
			assign ap_sbclr = ap[25];
			assign ap_sbinv = ap[24];
			assign ap_sbext = ap[23];
		end
		else begin
			assign ap_sbset = 1'b0;
			assign ap_sbclr = 1'b0;
			assign ap_sbinv = 1'b0;
			assign ap_sbext = 1'b0;
		end
	endgenerate
	generate
		if (pt[2187-:5] == 1) begin
			assign ap_slo = ap[38];
			assign ap_sro = ap[37];
		end
		else begin
			assign ap_slo = 1'b0;
			assign ap_sro = 1'b0;
		end
	endgenerate
	generate
		if (pt[2212-:5] == 1) begin
			assign ap_sh1add = ap[22];
			assign ap_sh2add = ap[21];
			assign ap_sh3add = ap[20];
			assign ap_zba = ap[19];
		end
		else begin
			assign ap_sh1add = 1'b0;
			assign ap_sh2add = 1'b0;
			assign ap_sh3add = 1'b0;
			assign ap_zba = 1'b0;
		end
	endgenerate
	rvdffpcie #(.WIDTH(31)) i_pc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(enable),
		.din(pc_in[31:1]),
		.dout(pc_ff[31:1])
	);
	rvdffe #(.WIDTH(32)) i_result_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(enable & valid_in),
		.din(result[31:0]),
		.dout(result_ff[31:0])
	);
	assign zba_a_in[31:0] = ((({32 {ap_sh1add}} & {a_in[30:0], 1'b0}) | ({32 {ap_sh2add}} & {a_in[29:0], 2'b00})) | ({32 {ap_sh3add}} & {a_in[28:0], 3'b000})) | ({32 {~ap_zba}} & a_in[31:0]);
	wire [31:0] bm;
	assign bm[31:0] = (ap[7] ? ~b_in[31:0] : b_in[31:0]);
	assign {cout, aout[31:0]} = ({1'b0, zba_a_in[31:0]} + {1'b0, bm[31:0]}) + {32'b00000000000000000000000000000000, ap[7]};
	assign ov = ((~a_in[31] & ~bm[31]) & aout[31]) | ((a_in[31] & bm[31]) & ~aout[31]);
	assign lt = (~ap[5] & (neg ^ ov)) | (ap[5] & ~cout);
	assign eq = a_in[31:0] == b_in[31:0];
	assign ne = ~eq;
	assign neg = aout[31];
	assign ge = ~lt;
	assign lout[31:0] = (((((({32 {csr_ren_in}} & csr_rddata_in[31:0]) | (({32 {ap[18] & ~ap_zbb}} & a_in[31:0]) & b_in[31:0])) | ({32 {ap[17] & ~ap_zbb}} & (a_in[31:0] | b_in[31:0]))) | ({32 {ap[16] & ~ap_zbb}} & (a_in[31:0] ^ b_in[31:0]))) | (({32 {ap[18] & ap_zbb}} & a_in[31:0]) & ~b_in[31:0])) | ({32 {ap[17] & ap_zbb}} & (a_in[31:0] | ~b_in[31:0]))) | ({32 {ap[16] & ap_zbb}} & (a_in[31:0] ^ ~b_in[31:0]));
	wire [5:0] shift_amount;
	wire [31:0] shift_mask;
	wire [62:0] shift_extend;
	wire [62:0] shift_long;
	assign shift_amount[5:0] = ((((((({6 {ap[15]}} & (6'd32 - {1'b0, b_in[4:0]})) | ({6 {ap[14]}} & {1'b0, b_in[4:0]})) | ({6 {ap[13]}} & {1'b0, b_in[4:0]})) | ({6 {ap_rol}} & (6'd32 - {1'b0, b_in[4:0]}))) | ({6 {ap_ror}} & {1'b0, b_in[4:0]})) | ({6 {ap_slo}} & (6'd32 - {1'b0, b_in[4:0]}))) | ({6 {ap_sro}} & {1'b0, b_in[4:0]})) | ({6 {ap_sbext}} & {1'b0, b_in[4:0]});
	assign shift_mask[31:0] = 32'hffffffff << ({5 {ap[15] | ap_slo}} & b_in[4:0]);
	assign shift_extend[31:0] = a_in[31:0];
	assign shift_extend[62:32] = ((((({31 {ap[13]}} & {31 {a_in[31]}}) | ({31 {ap[15]}} & a_in[30:0])) | ({31 {ap_rol}} & a_in[30:0])) | ({31 {ap_ror}} & a_in[30:0])) | ({31 {ap_slo}} & a_in[30:0])) | ({31 {ap_sro}} & {31 {1'b1}});
	assign shift_long[62:0] = shift_extend[62:0] >> shift_amount[4:0];
	assign sout[31:0] = (shift_long[31:0] & shift_mask[31:0]) | ({32 {ap_slo}} & ~shift_mask[31:0]);
	wire bitmanip_clz_ctz_sel;
	wire [31:0] bitmanip_a_reverse_ff;
	wire [31:0] bitmanip_lzd_in;
	reg [5:0] bitmanip_dw_lzd_enc;
	wire [5:0] bitmanip_clz_ctz_result;
	assign bitmanip_clz_ctz_sel = ap_clz | ap_ctz;
	assign bitmanip_a_reverse_ff[31:0] = {a_in[0], a_in[1], a_in[2], a_in[3], a_in[4], a_in[5], a_in[6], a_in[7], a_in[8], a_in[9], a_in[10], a_in[11], a_in[12], a_in[13], a_in[14], a_in[15], a_in[16], a_in[17], a_in[18], a_in[19], a_in[20], a_in[21], a_in[22], a_in[23], a_in[24], a_in[25], a_in[26], a_in[27], a_in[28], a_in[29], a_in[30], a_in[31]};
	assign bitmanip_lzd_in[31:0] = ({32 {ap_clz}} & a_in[31:0]) | ({32 {ap_ctz}} & bitmanip_a_reverse_ff[31:0]);
	reg [31:0] bitmanip_lzd_os;
	integer i;
	reg found;
	always @(*) begin
		bitmanip_lzd_os[31:0] = bitmanip_lzd_in[31:0];
		bitmanip_dw_lzd_enc[5:0] = 6'b000000;
		found = 1'b0;
		begin : sv2v_autoblock_42
			reg signed [31:0] i;
			for (i = 0; (i < 32) && (found == 0); i = i + 1)
				if (bitmanip_lzd_os[31] == 1'b0) begin
					bitmanip_dw_lzd_enc[5:0] = bitmanip_dw_lzd_enc[5:0] + 6'b000001;
					bitmanip_lzd_os[31:0] = bitmanip_lzd_os[31:0] << 1;
				end
				else
					found = 1'b1;
		end
	end
	assign bitmanip_clz_ctz_result[5:0] = {6 {bitmanip_clz_ctz_sel}} & {bitmanip_dw_lzd_enc[5], {5 {~bitmanip_dw_lzd_enc[5]}} & bitmanip_dw_lzd_enc[4:0]};
	reg [5:0] bitmanip_pcnt;
	wire [5:0] bitmanip_pcnt_result;
	integer bitmanip_pcnt_i;
	always @(*) begin
		bitmanip_pcnt[5:0] = 6'b000000;
		for (bitmanip_pcnt_i = 0; bitmanip_pcnt_i < 32; bitmanip_pcnt_i = bitmanip_pcnt_i + 1)
			bitmanip_pcnt[5:0] = bitmanip_pcnt[5:0] + {5'b00000, a_in[bitmanip_pcnt_i]};
	end
	assign bitmanip_pcnt_result[5:0] = {6 {ap_pcnt}} & bitmanip_pcnt[5:0];
	wire [31:0] bitmanip_sext_result;
	assign bitmanip_sext_result[31:0] = ({32 {ap_sext_b}} & {{24 {a_in[7]}}, a_in[7:0]}) | ({32 {ap_sext_h}} & {{16 {a_in[15]}}, a_in[15:0]});
	wire bitmanip_minmax_sel;
	wire [31:0] bitmanip_minmax_result;
	assign bitmanip_minmax_sel = ap_min | ap_max;
	wire bitmanip_minmax_sel_a;
	assign bitmanip_minmax_sel_a = ge ^ ap_min;
	assign bitmanip_minmax_result[31:0] = ({32 {bitmanip_minmax_sel & bitmanip_minmax_sel_a}} & a_in[31:0]) | ({32 {bitmanip_minmax_sel & ~bitmanip_minmax_sel_a}} & b_in[31:0]);
	wire [31:0] bitmanip_pack_result;
	wire [31:0] bitmanip_packu_result;
	wire [31:0] bitmanip_packh_result;
	assign bitmanip_pack_result[31:0] = {32 {ap_pack}} & {b_in[15:0], a_in[15:0]};
	assign bitmanip_packu_result[31:0] = {32 {ap_packu}} & {b_in[31:16], a_in[31:16]};
	assign bitmanip_packh_result[31:0] = {32 {ap_packh}} & {16'b0000000000000000, b_in[7:0], a_in[7:0]};
	wire [31:0] bitmanip_rev_result;
	wire [31:0] bitmanip_rev8_result;
	wire [31:0] bitmanip_orc_b_result;
	wire [31:0] bitmanip_orc16_result;
	assign bitmanip_rev_result[31:0] = {32 {ap_rev}} & {a_in[0], a_in[1], a_in[2], a_in[3], a_in[4], a_in[5], a_in[6], a_in[7], a_in[8], a_in[9], a_in[10], a_in[11], a_in[12], a_in[13], a_in[14], a_in[15], a_in[16], a_in[17], a_in[18], a_in[19], a_in[20], a_in[21], a_in[22], a_in[23], a_in[24], a_in[25], a_in[26], a_in[27], a_in[28], a_in[29], a_in[30], a_in[31]};
	assign bitmanip_rev8_result[31:0] = {32 {ap_rev8}} & {a_in[7:0], a_in[15:8], a_in[23:16], a_in[31:24]};
	assign bitmanip_orc_b_result[31:0] = {32 {ap_orc_b}} & {{8 {|a_in[31:24]}}, {8 {|a_in[23:16]}}, {8 {|a_in[15:8]}}, {8 {|a_in[7:0]}}};
	assign bitmanip_orc16_result[31:0] = {32 {ap_orc16}} & {{a_in[31:16] | a_in[15:0]}, {a_in[31:16] | a_in[15:0]}};
	wire [31:0] bitmanip_sb_1hot;
	wire [31:0] bitmanip_sb_data;
	assign bitmanip_sb_1hot[31:0] = 32'h00000001 << b_in[4:0];
	assign bitmanip_sb_data[31:0] = (({32 {ap_sbset}} & (a_in[31:0] | bitmanip_sb_1hot[31:0])) | ({32 {ap_sbclr}} & (a_in[31:0] & ~bitmanip_sb_1hot[31:0]))) | ({32 {ap_sbinv}} & (a_in[31:0] ^ bitmanip_sb_1hot[31:0]));
	assign sel_shift = (((((ap[15] | ap[14]) | ap[13]) | ap_slo) | ap_sro) | ap_rol) | ap_ror;
	assign sel_adder = ((((ap[8] | ap[7]) | ap_zba) & ~ap[6]) & ~ap_min) & ~ap_max;
	assign sel_pc = ((ap[4] | pp_in[34]) | pp_in[33]) | pp_in[31];
	assign csr_write_data[31:0] = (ap[0] ? b_in[31:0] : a_in[31:0]);
	assign slt_one = ap[6] & lt;
	assign result[31:0] = (((((((((((((((((lout[31:0] | ({32 {sel_shift}} & sout[31:0])) | ({32 {sel_adder}} & aout[31:0])) | ({32 {sel_pc}} & {pcout[31:1], 1'b0})) | ({32 {ap[1]}} & csr_write_data[31:0])) | {31'b0000000000000000000000000000000, slt_one}) | ({32 {ap_sbext}} & {31'b0000000000000000000000000000000, sout[0]})) | {26'b00000000000000000000000000, bitmanip_clz_ctz_result[5:0]}) | {26'b00000000000000000000000000, bitmanip_pcnt_result[5:0]}) | bitmanip_sext_result[31:0]) | bitmanip_minmax_result[31:0]) | bitmanip_pack_result[31:0]) | bitmanip_packu_result[31:0]) | bitmanip_packh_result[31:0]) | bitmanip_rev_result[31:0]) | bitmanip_rev8_result[31:0]) | bitmanip_orc_b_result[31:0]) | bitmanip_orc16_result[31:0]) | bitmanip_sb_data[31:0];
	assign any_jal = ((ap[4] | pp_in[34]) | pp_in[33]) | pp_in[31];
	assign actual_taken = ((((ap[12] & eq) | (ap[11] & ne)) | (ap[10] & lt)) | (ap[9] & ge)) | any_jal;
	rvbradder ibradder(
		.pc(pc_in[31:1]),
		.offset(brimm_in[12:1]),
		.dout(pcout[31:1])
	);
	assign pred_correct_out = (((valid_in & ap[2]) & ~actual_taken) & ~any_jal) | (((valid_in & ap[3]) & actual_taken) & ~any_jal);
	assign flush_path_out[31:1] = (any_jal ? aout[31:1] : pcout[31:1]);
	assign cond_mispredict = (ap[3] & ~actual_taken) | (ap[2] & actual_taken);
	assign target_mispredict = pp_in[31] & (pp_in[30:0] != aout[31:1]);
	assign flush_upper_out = ((((ap[4] | cond_mispredict) | target_mispredict) & valid_in) & ~flush_upper_x) & ~flush_lower_r;
	assign flush_final_out = ((((ap[4] | cond_mispredict) | target_mispredict) & valid_in) & ~flush_upper_x) | flush_lower_r;
	assign newhist[1] = (pp_in[51] & pp_in[50]) | (~pp_in[50] & actual_taken);
	assign newhist[0] = (~pp_in[51] & ~actual_taken) | (pp_in[51] & actual_taken);
	always @(*) begin
		predict_p_out = pp_in;
		predict_p_out[55] = (~flush_upper_x & ~flush_lower_r) & (cond_mispredict | target_mispredict);
		predict_p_out[54] = actual_taken;
		predict_p_out[51] = newhist[1];
		predict_p_out[50] = newhist[0];
	end
endmodule
module eb1_exu_div_ctl (
	clk,
	rst_l,
	scan_mode,
	dp,
	dividend,
	divisor,
	cancel,
	finish_dly,
	out
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire [2:0] dp;
	input wire [31:0] dividend;
	input wire [31:0] divisor;
	input wire cancel;
	output wire finish_dly;
	output wire [31:0] out;
	wire [31:0] out_raw;
	assign out[31:0] = {32 {finish_dly}} & out_raw[31:0];
	generate
		if (pt[1262-:5] == 0) eb1_exu_div_existing_1bit_cheapshortq i_existing_1bit_div_cheapshortq(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.cancel(cancel),
			.valid_in(dp[2]),
			.signed_in(~dp[1]),
			.rem_in(dp[0]),
			.dividend_in(dividend[31:0]),
			.divisor_in(divisor[31:0]),
			.valid_out(finish_dly),
			.data_out(out_raw[31:0])
		);
	endgenerate
	generate
		if ((pt[1262-:5] == 1) & (pt[1269-:7] == 1)) eb1_exu_div_new_1bit_fullshortq i_new_1bit_div_fullshortq(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.cancel(cancel),
			.valid_in(dp[2]),
			.signed_in(~dp[1]),
			.rem_in(dp[0]),
			.dividend_in(dividend[31:0]),
			.divisor_in(divisor[31:0]),
			.valid_out(finish_dly),
			.data_out(out_raw[31:0])
		);
	endgenerate
	generate
		if ((pt[1262-:5] == 1) & (pt[1269-:7] == 2)) eb1_exu_div_new_2bit_fullshortq i_new_2bit_div_fullshortq(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.cancel(cancel),
			.valid_in(dp[2]),
			.signed_in(~dp[1]),
			.rem_in(dp[0]),
			.dividend_in(dividend[31:0]),
			.divisor_in(divisor[31:0]),
			.valid_out(finish_dly),
			.data_out(out_raw[31:0])
		);
	endgenerate
	generate
		if ((pt[1262-:5] == 1) & (pt[1269-:7] == 3)) eb1_exu_div_new_3bit_fullshortq i_new_3bit_div_fullshortq(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.cancel(cancel),
			.valid_in(dp[2]),
			.signed_in(~dp[1]),
			.rem_in(dp[0]),
			.dividend_in(dividend[31:0]),
			.divisor_in(divisor[31:0]),
			.valid_out(finish_dly),
			.data_out(out_raw[31:0])
		);
	endgenerate
	generate
		if ((pt[1262-:5] == 1) & (pt[1269-:7] == 4)) eb1_exu_div_new_4bit_fullshortq i_new_4bit_div_fullshortq(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.cancel(cancel),
			.valid_in(dp[2]),
			.signed_in(~dp[1]),
			.rem_in(dp[0]),
			.dividend_in(dividend[31:0]),
			.divisor_in(divisor[31:0]),
			.valid_out(finish_dly),
			.data_out(out_raw[31:0])
		);
	endgenerate
endmodule
module eb1_exu_div_existing_1bit_cheapshortq (
	clk,
	rst_l,
	scan_mode,
	cancel,
	valid_in,
	signed_in,
	rem_in,
	dividend_in,
	divisor_in,
	valid_out,
	data_out
);
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire cancel;
	input wire valid_in;
	input wire signed_in;
	input wire rem_in;
	input wire [31:0] dividend_in;
	input wire [31:0] divisor_in;
	output wire valid_out;
	output wire [31:0] data_out;
	wire div_clken;
	wire run_in;
	wire run_state;
	wire [5:0] count_in;
	wire [5:0] count;
	wire [32:0] m_ff;
	wire qff_enable;
	wire aff_enable;
	wire [32:0] q_in;
	wire [32:0] q_ff;
	wire [32:0] a_in;
	wire [32:0] a_ff;
	wire [32:0] m_eff;
	wire [32:0] a_shift;
	wire dividend_neg_ff;
	wire divisor_neg_ff;
	wire [31:0] dividend_comp;
	wire [31:0] dividend_eff;
	wire [31:0] q_ff_comp;
	wire [31:0] q_ff_eff;
	wire [31:0] a_ff_comp;
	wire [31:0] a_ff_eff;
	wire sign_ff;
	wire sign_eff;
	wire rem_ff;
	wire add;
	wire [32:0] a_eff;
	wire [64:0] a_eff_shift;
	wire rem_correct;
	wire valid_ff_x;
	wire valid_x;
	wire finish;
	wire finish_ff;
	wire smallnum_case;
	wire smallnum_case_ff;
	wire [3:0] smallnum;
	wire [3:0] smallnum_ff;
	wire m_already_comp;
	wire [4:0] a_cls;
	wire [4:0] b_cls;
	wire [5:0] shortq_shift;
	wire [5:0] shortq_shift_ff;
	wire [5:0] shortq;
	wire shortq_enable;
	wire shortq_enable_ff;
	wire [32:0] short_dividend;
	wire [3:0] shortq_raw;
	wire [3:0] shortq_shift_xx;
	rvdffe #(.WIDTH(23)) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(div_clken),
		.din({valid_in & ~cancel, finish & ~cancel, run_in, count_in[5:0], (valid_in & dividend_in[31]) | (~valid_in & dividend_neg_ff), (valid_in & divisor_in[31]) | (~valid_in & divisor_neg_ff), (valid_in & sign_eff) | (~valid_in & sign_ff), (valid_in & rem_in) | (~valid_in & rem_ff), smallnum_case, smallnum[3:0], shortq_enable, shortq_shift[3:0]}),
		.dout({valid_ff_x, finish_ff, run_state, count[5:0], dividend_neg_ff, divisor_neg_ff, sign_ff, rem_ff, smallnum_case_ff, smallnum_ff[3:0], shortq_enable_ff, shortq_shift_xx[3:0]})
	);
	rvdffe #(.WIDTH(33)) mff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(valid_in),
		.din({signed_in & divisor_in[31], divisor_in[31:0]}),
		.dout(m_ff[32:0])
	);
	rvdffe #(.WIDTH(33)) qff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qff_enable),
		.din(q_in[32:0]),
		.dout(q_ff[32:0])
	);
	rvdffe #(.WIDTH(33)) aff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(aff_enable),
		.din(a_in[32:0]),
		.dout(a_ff[32:0])
	);
	rvtwoscomp #(.WIDTH(32)) i_dividend_comp(
		.din(q_ff[31:0]),
		.dout(dividend_comp[31:0])
	);
	rvtwoscomp #(.WIDTH(32)) i_q_ff_comp(
		.din(q_ff[31:0]),
		.dout(q_ff_comp[31:0])
	);
	rvtwoscomp #(.WIDTH(32)) i_a_ff_comp(
		.din(a_ff[31:0]),
		.dout(a_ff_comp[31:0])
	);
	assign valid_x = valid_ff_x & ~cancel;
	assign smallnum_case = (((((q_ff[31:4] == 28'b0000000000000000000000000000) & (m_ff[31:4] == 28'b0000000000000000000000000000)) & (m_ff[31:0] != 32'b00000000000000000000000000000000)) & ~rem_ff) & valid_x) | ((((q_ff[31:0] == 32'b00000000000000000000000000000000) & (m_ff[31:0] != 32'b00000000000000000000000000000000)) & ~rem_ff) & valid_x);
	assign smallnum[3] = ((q_ff[3] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[1];
	assign smallnum[2] = ((((q_ff[3] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[0]) | (((q_ff[2] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[1])) | (((q_ff[3] & q_ff[2]) & ~m_ff[3]) & ~m_ff[2]);
	assign smallnum[1] = ((((((((((q_ff[2] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[0]) | (((q_ff[1] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[1])) | (((q_ff[3] & ~m_ff[3]) & ~m_ff[1]) & ~m_ff[0])) | (((((q_ff[3] & ~q_ff[2]) & ~m_ff[3]) & ~m_ff[2]) & m_ff[1]) & m_ff[0])) | ((((~q_ff[3] & q_ff[2]) & q_ff[1]) & ~m_ff[3]) & ~m_ff[2])) | (((q_ff[3] & q_ff[2]) & ~m_ff[3]) & ~m_ff[0])) | ((((q_ff[3] & q_ff[2]) & ~m_ff[3]) & m_ff[2]) & ~m_ff[1])) | (((q_ff[3] & q_ff[1]) & ~m_ff[3]) & ~m_ff[1])) | ((((q_ff[3] & q_ff[2]) & q_ff[1]) & ~m_ff[3]) & m_ff[2]);
	assign smallnum[0] = ((((((((((((((((((((((((((((q_ff[2] & q_ff[1]) & q_ff[0]) & ~m_ff[3]) & ~m_ff[1]) | (((((q_ff[3] & ~q_ff[2]) & q_ff[0]) & ~m_ff[3]) & m_ff[1]) & m_ff[0])) | (((q_ff[2] & ~m_ff[3]) & ~m_ff[1]) & ~m_ff[0])) | (((q_ff[1] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[0])) | (((q_ff[0] & ~m_ff[3]) & ~m_ff[2]) & ~m_ff[1])) | ((((((~q_ff[3] & q_ff[2]) & ~q_ff[1]) & ~m_ff[3]) & ~m_ff[2]) & m_ff[1]) & m_ff[0])) | ((((~q_ff[3] & q_ff[2]) & q_ff[1]) & ~m_ff[3]) & ~m_ff[0])) | (((q_ff[3] & ~m_ff[2]) & ~m_ff[1]) & ~m_ff[0])) | ((((q_ff[3] & ~q_ff[2]) & ~m_ff[3]) & m_ff[2]) & m_ff[1])) | (((((~q_ff[3] & q_ff[2]) & q_ff[1]) & ~m_ff[3]) & m_ff[2]) & ~m_ff[1])) | ((((~q_ff[3] & q_ff[2]) & q_ff[0]) & ~m_ff[3]) & ~m_ff[1])) | (((((q_ff[3] & ~q_ff[2]) & ~q_ff[1]) & ~m_ff[3]) & m_ff[2]) & m_ff[0])) | ((((~q_ff[2] & q_ff[1]) & q_ff[0]) & ~m_ff[3]) & ~m_ff[2])) | (((q_ff[3] & q_ff[2]) & ~m_ff[1]) & ~m_ff[0])) | (((q_ff[3] & q_ff[1]) & ~m_ff[2]) & ~m_ff[0])) | (((((~q_ff[3] & q_ff[2]) & q_ff[1]) & q_ff[0]) & ~m_ff[3]) & m_ff[2])) | (((q_ff[3] & q_ff[2]) & m_ff[3]) & ~m_ff[2])) | ((((q_ff[3] & q_ff[1]) & m_ff[3]) & ~m_ff[2]) & ~m_ff[1])) | (((q_ff[3] & q_ff[0]) & ~m_ff[2]) & ~m_ff[1])) | (((((q_ff[3] & ~q_ff[1]) & ~m_ff[3]) & m_ff[2]) & m_ff[1]) & m_ff[0])) | ((((q_ff[3] & q_ff[2]) & q_ff[1]) & m_ff[3]) & ~m_ff[0])) | ((((q_ff[3] & q_ff[2]) & q_ff[1]) & m_ff[3]) & ~m_ff[1])) | ((((q_ff[3] & q_ff[2]) & q_ff[0]) & m_ff[3]) & ~m_ff[1])) | ((((q_ff[3] & ~q_ff[2]) & q_ff[1]) & ~m_ff[3]) & m_ff[1])) | (((q_ff[3] & q_ff[1]) & q_ff[0]) & ~m_ff[2])) | ((((q_ff[3] & q_ff[2]) & q_ff[1]) & q_ff[0]) & m_ff[3]);
	assign short_dividend[31:0] = q_ff[31:0];
	assign short_dividend[32] = sign_ff & q_ff[31];
	assign a_cls[4:3] = 2'b00;
	assign a_cls[2] = (~short_dividend[32] & (short_dividend[31:24] != {8 {1'b0}})) | (short_dividend[32] & (short_dividend[31:23] != {9 {1'b1}}));
	assign a_cls[1] = (~short_dividend[32] & (short_dividend[23:16] != {8 {1'b0}})) | (short_dividend[32] & (short_dividend[22:15] != {8 {1'b1}}));
	assign a_cls[0] = (~short_dividend[32] & (short_dividend[15:8] != {8 {1'b0}})) | (short_dividend[32] & (short_dividend[14:7] != {8 {1'b1}}));
	assign b_cls[4:3] = 2'b00;
	assign b_cls[2] = (~m_ff[32] & (m_ff[31:24] != {8 {1'b0}})) | (m_ff[32] & (m_ff[31:24] != {8 {1'b1}}));
	assign b_cls[1] = (~m_ff[32] & (m_ff[23:16] != {8 {1'b0}})) | (m_ff[32] & (m_ff[23:16] != {8 {1'b1}}));
	assign b_cls[0] = (~m_ff[32] & (m_ff[15:8] != {8 {1'b0}})) | (m_ff[32] & (m_ff[15:8] != {8 {1'b1}}));
	assign shortq_raw[3] = ((((((a_cls[2:1] == 2'b01) & (b_cls[2] == 1'b1)) | ((a_cls[2:0] == 3'b001) & (b_cls[2] == 1'b1))) | ((a_cls[2:0] == 3'b000) & (b_cls[2] == 1'b1))) | ((a_cls[2:0] == 3'b001) & (b_cls[2:1] == 2'b01))) | ((a_cls[2:0] == 3'b000) & (b_cls[2:1] == 2'b01))) | ((a_cls[2:0] == 3'b000) & (b_cls[2:0] == 3'b001));
	assign shortq_raw[2] = ((((a_cls[2] == 1'b1) & (b_cls[2] == 1'b1)) | ((a_cls[2:1] == 2'b01) & (b_cls[2:1] == 2'b01))) | ((a_cls[2:0] == 3'b001) & (b_cls[2:0] == 3'b001))) | ((a_cls[2:0] == 3'b000) & (b_cls[2:0] == 3'b000));
	assign shortq_raw[1] = (((a_cls[2] == 1'b1) & (b_cls[2:1] == 2'b01)) | ((a_cls[2:1] == 2'b01) & (b_cls[2:0] == 3'b001))) | ((a_cls[2:0] == 3'b001) & (b_cls[2:0] == 3'b000));
	assign shortq_raw[0] = ((a_cls[2] == 1'b1) & (b_cls[2:0] == 3'b001)) | ((a_cls[2:1] == 2'b01) & (b_cls[2:0] == 3'b000));
	assign shortq_enable = (valid_ff_x & (m_ff[31:0] != 32'b00000000000000000000000000000000)) & (shortq_raw[3:0] != 4'b0000);
	assign shortq_shift[3:0] = {4 {shortq_enable}} & shortq_raw[3:0];
	assign shortq[5:0] = 6'b000000;
	assign shortq_shift[5:4] = 2'b00;
	assign shortq_shift_ff[5] = 1'b0;
	assign shortq_shift_ff[4:0] = ((({5 {shortq_shift_xx[3]}} & 5'b11111) | ({5 {shortq_shift_xx[2]}} & 5'b11000)) | ({5 {shortq_shift_xx[1]}} & 5'b10000)) | ({5 {shortq_shift_xx[0]}} & 5'b01000);
	assign div_clken = ((valid_in | run_state) | finish) | finish_ff;
	assign run_in = ((valid_in | run_state) & ~finish) & ~cancel;
	assign count_in[5:0] = {6 {((run_state & ~finish) & ~cancel) & ~shortq_enable}} & ((count[5:0] + {1'b0, shortq_shift_ff[4:0]}) + 6'd1);
	assign finish = smallnum_case | (~rem_ff ? count[5:0] == 6'd32 : count[5:0] == 6'd33);
	assign valid_out = finish_ff & ~cancel;
	assign sign_eff = signed_in & (divisor_in[31:0] != 32'b00000000000000000000000000000000);
	assign q_in[32:0] = (({33 {~run_state}} & {1'b0, dividend_in[31:0]}) | ({33 {run_state & (valid_ff_x | shortq_enable_ff)}} & ({dividend_eff[31:0], ~a_in[32]} << shortq_shift_ff[4:0]))) | ({33 {run_state & ~(valid_ff_x | shortq_enable_ff)}} & {q_ff[31:0], ~a_in[32]});
	assign qff_enable = valid_in | (run_state & ~shortq_enable);
	assign dividend_eff[31:0] = (sign_ff & dividend_neg_ff ? dividend_comp[31:0] : q_ff[31:0]);
	assign m_eff[32:0] = (add ? m_ff[32:0] : ~m_ff[32:0]);
	assign a_eff_shift[64:0] = {33'b000000000000000000000000000000000, dividend_eff[31:0]} << shortq_shift_ff[4:0];
	assign a_eff[32:0] = (({33 {rem_correct}} & a_ff[32:0]) | ({33 {~rem_correct & ~shortq_enable_ff}} & {a_ff[31:0], q_ff[32]})) | ({33 {~rem_correct & shortq_enable_ff}} & a_eff_shift[64:32]);
	assign a_shift[32:0] = {33 {run_state}} & a_eff[32:0];
	assign a_in[32:0] = {33 {run_state}} & ((a_shift[32:0] + m_eff[32:0]) + {32'b00000000000000000000000000000000, ~add});
	assign aff_enable = (valid_in | ((run_state & ~shortq_enable) & (count[5:0] != 6'd33))) | rem_correct;
	assign m_already_comp = divisor_neg_ff & sign_ff;
	assign add = (a_ff[32] | rem_correct) ^ m_already_comp;
	assign rem_correct = ((count[5:0] == 6'd33) & rem_ff) & a_ff[32];
	assign q_ff_eff[31:0] = (sign_ff & (dividend_neg_ff ^ divisor_neg_ff) ? q_ff_comp[31:0] : q_ff[31:0]);
	assign a_ff_eff[31:0] = (sign_ff & dividend_neg_ff ? a_ff_comp[31:0] : a_ff[31:0]);
	assign data_out[31:0] = (({32 {smallnum_case_ff}} & {28'b0000000000000000000000000000, smallnum_ff[3:0]}) | ({32 {rem_ff}} & a_ff_eff[31:0])) | ({32 {~smallnum_case_ff & ~rem_ff}} & q_ff_eff[31:0]);
endmodule
module eb1_exu_div_new_1bit_fullshortq (
	clk,
	rst_l,
	scan_mode,
	cancel,
	valid_in,
	signed_in,
	rem_in,
	dividend_in,
	divisor_in,
	valid_out,
	data_out
);
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire cancel;
	input wire valid_in;
	input wire signed_in;
	input wire rem_in;
	input wire [31:0] dividend_in;
	input wire [31:0] divisor_in;
	output wire valid_out;
	output wire [31:0] data_out;
	wire valid_ff_in;
	wire valid_ff;
	wire finish_raw;
	wire finish;
	wire finish_ff;
	wire running_state;
	wire misc_enable;
	wire [2:0] control_in;
	wire [2:0] control_ff;
	wire dividend_sign_ff;
	wire divisor_sign_ff;
	wire rem_ff;
	wire count_enable;
	wire [6:0] count_in;
	wire [6:0] count_ff;
	wire smallnum_case;
	wire [3:0] smallnum;
	wire a_enable;
	wire a_shift;
	wire [31:0] a_in;
	wire [31:0] a_ff;
	wire b_enable;
	wire b_twos_comp;
	wire [32:0] b_in;
	wire [32:0] b_ff;
	wire [31:0] q_in;
	wire [31:0] q_ff;
	wire rq_enable;
	wire r_sign_sel;
	wire r_restore_sel;
	wire r_adder_sel;
	wire [31:0] r_in;
	wire [31:0] r_ff;
	wire twos_comp_q_sel;
	wire twos_comp_b_sel;
	wire [31:0] twos_comp_in;
	wire [31:0] twos_comp_out;
	wire quotient_set;
	wire [32:0] adder_out;
	wire [63:0] ar_shifted;
	wire [5:0] shortq;
	wire [4:0] shortq_shift;
	wire [4:0] shortq_shift_ff;
	wire shortq_enable;
	wire shortq_enable_ff;
	wire [32:0] shortq_dividend;
	wire by_zero_case;
	wire by_zero_case_ff;
	rvdffe #(.WIDTH(19)) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(misc_enable),
		.din({valid_ff_in, control_in[2:0], by_zero_case, shortq_enable, shortq_shift[4:0], finish, count_in[6:0]}),
		.dout({valid_ff, control_ff[2:0], by_zero_case_ff, shortq_enable_ff, shortq_shift_ff[4:0], finish_ff, count_ff[6:0]})
	);
	rvdffe #(.WIDTH(32)) i_a_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(a_enable),
		.din(a_in[31:0]),
		.dout(a_ff[31:0])
	);
	rvdffe #(.WIDTH(33)) i_b_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(b_enable),
		.din(b_in[32:0]),
		.dout(b_ff[32:0])
	);
	rvdffe #(.WIDTH(32)) i_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(r_in[31:0]),
		.dout(r_ff[31:0])
	);
	rvdffe #(.WIDTH(32)) i_q_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(q_in[31:0]),
		.dout(q_ff[31:0])
	);
	assign valid_ff_in = valid_in & ~cancel;
	assign control_in[2] = (~valid_in & control_ff[2]) | ((valid_in & signed_in) & dividend_in[31]);
	assign control_in[1] = (~valid_in & control_ff[1]) | ((valid_in & signed_in) & divisor_in[31]);
	assign control_in[0] = (~valid_in & control_ff[0]) | (valid_in & rem_in);
	assign dividend_sign_ff = control_ff[2];
	assign divisor_sign_ff = control_ff[1];
	assign rem_ff = control_ff[0];
	assign by_zero_case = valid_ff & (b_ff[31:0] == 32'b00000000000000000000000000000000);
	assign misc_enable = (((valid_in | valid_ff) | cancel) | running_state) | finish_ff;
	assign running_state = |count_ff[6:0] | shortq_enable_ff;
	assign finish_raw = (smallnum_case | by_zero_case) | (count_ff[6:0] == 7'd32);
	assign finish = finish_raw & ~cancel;
	assign count_enable = ((((valid_ff | running_state) & ~finish) & ~finish_ff) & ~cancel) & ~shortq_enable;
	assign count_in[6:0] = {7 {count_enable}} & ((count_ff[6:0] + 7'b0000001) + {2'b00, shortq_shift_ff[4:0]});
	assign a_enable = valid_in | running_state;
	assign a_shift = running_state & ~shortq_enable_ff;
	assign ar_shifted[63:0] = {{32 {dividend_sign_ff}}, a_ff[31:0]} << shortq_shift_ff[4:0];
	assign a_in[31:0] = (({32 {~a_shift & ~shortq_enable_ff}} & dividend_in[31:0]) | ({32 {a_shift}} & {a_ff[30:0], 1'b0})) | ({32 {shortq_enable_ff}} & ar_shifted[31:0]);
	assign b_enable = valid_in | b_twos_comp;
	assign b_twos_comp = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign b_in[32:0] = ({33 {~b_twos_comp}} & {signed_in & divisor_in[31], divisor_in[31:0]}) | ({33 {b_twos_comp}} & {~divisor_sign_ff, twos_comp_out[31:0]});
	assign rq_enable = (valid_in | valid_ff) | running_state;
	assign r_sign_sel = (valid_ff & dividend_sign_ff) & ~by_zero_case;
	assign r_restore_sel = (running_state & ~quotient_set) & ~shortq_enable_ff;
	assign r_adder_sel = (running_state & quotient_set) & ~shortq_enable_ff;
	assign r_in[31:0] = (((({32 {r_sign_sel}} & 32'hffffffff) | ({32 {r_restore_sel}} & {r_ff[30:0], a_ff[31]})) | ({32 {r_adder_sel}} & adder_out[31:0])) | ({32 {shortq_enable_ff}} & ar_shifted[63:32])) | ({32 {by_zero_case}} & a_ff[31:0]);
	assign q_in[31:0] = (({32 {~valid_ff}} & {q_ff[30:0], quotient_set}) | ({32 {smallnum_case}} & {28'b0000000000000000000000000000, smallnum[3:0]})) | ({32 {by_zero_case}} & {32 {1'b1}});
	assign adder_out[32:0] = {r_ff[31:0], a_ff[31]} + {b_ff[32:0]};
	assign quotient_set = (~adder_out[32] ^ dividend_sign_ff) | ((a_ff[30:0] == 31'b0000000000000000000000000000000) & (adder_out[32:0] == 33'b000000000000000000000000000000000));
	assign twos_comp_b_sel = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign twos_comp_q_sel = ((~valid_ff & ~rem_ff) & (dividend_sign_ff ^ divisor_sign_ff)) & ~by_zero_case_ff;
	assign twos_comp_in[31:0] = ({32 {twos_comp_q_sel}} & q_ff[31:0]) | ({32 {twos_comp_b_sel}} & b_ff[31:0]);
	rvtwoscomp #(.WIDTH(32)) i_twos_comp(
		.din(twos_comp_in[31:0]),
		.dout(twos_comp_out[31:0])
	);
	assign valid_out = finish_ff & ~cancel;
	assign data_out[31:0] = (({32 {~rem_ff & ~twos_comp_q_sel}} & q_ff[31:0]) | ({32 {rem_ff}} & r_ff[31:0])) | ({32 {twos_comp_q_sel}} & twos_comp_out[31:0]);
	assign smallnum_case = ((((((a_ff[31:4] == 28'b0000000000000000000000000000) & (b_ff[31:4] == 28'b0000000000000000000000000000)) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel) | (((((a_ff[31:0] == 32'b00000000000000000000000000000000) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel);
	assign smallnum[3] = ((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1];
	assign smallnum[2] = ((((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[2]);
	assign smallnum[1] = ((((((((((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[1]) & ~b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]);
	assign smallnum[0] = ((((((((((((((((((((((((((((a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1]) | (((((a_ff[3] & ~a_ff[2]) & a_ff[0]) & ~b_ff[3]) & b_ff[1]) & b_ff[0])) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0])) | (((a_ff[0] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | ((((((~a_ff[3] & a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[0])) | (((a_ff[3] & ~b_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | ((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & b_ff[2]) & b_ff[1])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | ((((~a_ff[3] & a_ff[2]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[0])) | ((((~a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[3] & a_ff[1]) & ~b_ff[2]) & ~b_ff[0])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & b_ff[2])) | (((a_ff[3] & a_ff[2]) & b_ff[3]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[1]) & b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[0]) & ~b_ff[2]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[0]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & ~a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[1])) | (((a_ff[3] & a_ff[1]) & a_ff[0]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & b_ff[3]);
	assign shortq_dividend[32:0] = {dividend_sign_ff, a_ff[31:0]};
	wire [5:0] dw_a_enc;
	wire [5:0] dw_b_enc;
	wire [6:0] dw_shortq_raw;
	eb1_exu_div_cls i_a_cls(
		.operand(shortq_dividend[32:0]),
		.cls(dw_a_enc[4:0])
	);
	eb1_exu_div_cls i_b_cls(
		.operand(b_ff[32:0]),
		.cls(dw_b_enc[4:0])
	);
	assign dw_a_enc[5] = 1'b0;
	assign dw_b_enc[5] = 1'b0;
	assign dw_shortq_raw[6:0] = ({1'b0, dw_b_enc[5:0]} - {1'b0, dw_a_enc[5:0]}) + 7'd1;
	assign shortq[5:0] = (dw_shortq_raw[6] ? 6'd0 : dw_shortq_raw[5:0]);
	assign shortq_enable = ((valid_ff & ~shortq[5]) & ~(shortq[4:1] == 4'b1111)) & ~cancel;
	assign shortq_shift[4:0] = (~shortq_enable ? 5'd0 : 5'b11111 - shortq[4:0]);
endmodule
module eb1_exu_div_new_2bit_fullshortq (
	clk,
	rst_l,
	scan_mode,
	cancel,
	valid_in,
	signed_in,
	rem_in,
	dividend_in,
	divisor_in,
	valid_out,
	data_out
);
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire cancel;
	input wire valid_in;
	input wire signed_in;
	input wire rem_in;
	input wire [31:0] dividend_in;
	input wire [31:0] divisor_in;
	output wire valid_out;
	output wire [31:0] data_out;
	wire valid_ff_in;
	wire valid_ff;
	wire finish_raw;
	wire finish;
	wire finish_ff;
	wire running_state;
	wire misc_enable;
	wire [2:0] control_in;
	wire [2:0] control_ff;
	wire dividend_sign_ff;
	wire divisor_sign_ff;
	wire rem_ff;
	wire count_enable;
	wire [6:0] count_in;
	wire [6:0] count_ff;
	wire smallnum_case;
	wire [3:0] smallnum;
	wire a_enable;
	wire a_shift;
	wire [31:0] a_in;
	wire [31:0] a_ff;
	wire b_enable;
	wire b_twos_comp;
	wire [32:0] b_in;
	wire [34:0] b_ff;
	wire [31:0] q_in;
	wire [31:0] q_ff;
	wire rq_enable;
	wire r_sign_sel;
	wire r_restore_sel;
	wire r_adder1_sel;
	wire r_adder2_sel;
	wire r_adder3_sel;
	wire [31:0] r_in;
	wire [31:0] r_ff;
	wire twos_comp_q_sel;
	wire twos_comp_b_sel;
	wire [31:0] twos_comp_in;
	wire [31:0] twos_comp_out;
	wire [3:1] quotient_raw;
	wire [1:0] quotient_new;
	wire [32:0] adder1_out;
	wire [33:0] adder2_out;
	wire [34:0] adder3_out;
	wire [63:0] ar_shifted;
	wire [5:0] shortq;
	wire [4:0] shortq_shift;
	wire [4:1] shortq_shift_ff;
	wire shortq_enable;
	wire shortq_enable_ff;
	wire [32:0] shortq_dividend;
	wire by_zero_case;
	wire by_zero_case_ff;
	rvdffe #(.WIDTH(18)) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(misc_enable),
		.din({valid_ff_in, control_in[2:0], by_zero_case, shortq_enable, shortq_shift[4:1], finish, count_in[6:0]}),
		.dout({valid_ff, control_ff[2:0], by_zero_case_ff, shortq_enable_ff, shortq_shift_ff[4:1], finish_ff, count_ff[6:0]})
	);
	rvdffe #(.WIDTH(32)) i_a_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(a_enable),
		.din(a_in[31:0]),
		.dout(a_ff[31:0])
	);
	rvdffe #(.WIDTH(33)) i_b_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(b_enable),
		.din(b_in[32:0]),
		.dout(b_ff[32:0])
	);
	rvdffe #(.WIDTH(32)) i_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(r_in[31:0]),
		.dout(r_ff[31:0])
	);
	rvdffe #(.WIDTH(32)) i_q_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(q_in[31:0]),
		.dout(q_ff[31:0])
	);
	assign valid_ff_in = valid_in & ~cancel;
	assign control_in[2] = (~valid_in & control_ff[2]) | ((valid_in & signed_in) & dividend_in[31]);
	assign control_in[1] = (~valid_in & control_ff[1]) | ((valid_in & signed_in) & divisor_in[31]);
	assign control_in[0] = (~valid_in & control_ff[0]) | (valid_in & rem_in);
	assign dividend_sign_ff = control_ff[2];
	assign divisor_sign_ff = control_ff[1];
	assign rem_ff = control_ff[0];
	assign by_zero_case = valid_ff & (b_ff[31:0] == 32'b00000000000000000000000000000000);
	assign misc_enable = (((valid_in | valid_ff) | cancel) | running_state) | finish_ff;
	assign running_state = |count_ff[6:0] | shortq_enable_ff;
	assign finish_raw = (smallnum_case | by_zero_case) | (count_ff[6:0] == 7'd32);
	assign finish = finish_raw & ~cancel;
	assign count_enable = ((((valid_ff | running_state) & ~finish) & ~finish_ff) & ~cancel) & ~shortq_enable;
	assign count_in[6:0] = {7 {count_enable}} & ((count_ff[6:0] + 7'b0000010) + {2'b00, shortq_shift_ff[4:1], 1'b0});
	assign a_enable = valid_in | running_state;
	assign a_shift = running_state & ~shortq_enable_ff;
	assign ar_shifted[63:0] = {{32 {dividend_sign_ff}}, a_ff[31:0]} << {shortq_shift_ff[4:1], 1'b0};
	assign a_in[31:0] = (({32 {~a_shift & ~shortq_enable_ff}} & dividend_in[31:0]) | ({32 {a_shift}} & {a_ff[29:0], 2'b00})) | ({32 {shortq_enable_ff}} & ar_shifted[31:0]);
	assign b_enable = valid_in | b_twos_comp;
	assign b_twos_comp = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign b_in[32:0] = ({33 {~b_twos_comp}} & {signed_in & divisor_in[31], divisor_in[31:0]}) | ({33 {b_twos_comp}} & {~divisor_sign_ff, twos_comp_out[31:0]});
	assign rq_enable = (valid_in | valid_ff) | running_state;
	assign r_sign_sel = (valid_ff & dividend_sign_ff) & ~by_zero_case;
	assign r_restore_sel = (running_state & (quotient_new[1:0] == 2'b00)) & ~shortq_enable_ff;
	assign r_adder1_sel = (running_state & (quotient_new[1:0] == 2'b01)) & ~shortq_enable_ff;
	assign r_adder2_sel = (running_state & (quotient_new[1:0] == 2'b10)) & ~shortq_enable_ff;
	assign r_adder3_sel = (running_state & (quotient_new[1:0] == 2'b11)) & ~shortq_enable_ff;
	assign r_in[31:0] = (((((({32 {r_sign_sel}} & 32'hffffffff) | ({32 {r_restore_sel}} & {r_ff[29:0], a_ff[31:30]})) | ({32 {r_adder1_sel}} & adder1_out[31:0])) | ({32 {r_adder2_sel}} & adder2_out[31:0])) | ({32 {r_adder3_sel}} & adder3_out[31:0])) | ({32 {shortq_enable_ff}} & ar_shifted[63:32])) | ({32 {by_zero_case}} & a_ff[31:0]);
	assign q_in[31:0] = (({32 {~valid_ff}} & {q_ff[29:0], quotient_new[1:0]}) | ({32 {smallnum_case}} & {28'b0000000000000000000000000000, smallnum[3:0]})) | ({32 {by_zero_case}} & {32 {1'b1}});
	assign b_ff[34:33] = {b_ff[32], b_ff[32]};
	assign adder1_out[32:0] = {r_ff[30:0], a_ff[31:30]} + b_ff[32:0];
	assign adder2_out[33:0] = {r_ff[31:0], a_ff[31:30]} + {b_ff[32:0], 1'b0};
	assign adder3_out[34:0] = ({r_ff[31], r_ff[31:0], a_ff[31:30]} + {b_ff[33:0], 1'b0}) + b_ff[34:0];
	assign quotient_raw[1] = (~adder1_out[32] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder1_out[32:0] == 33'b000000000000000000000000000000000));
	assign quotient_raw[2] = (~adder2_out[33] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder2_out[33:0] == 34'b0000000000000000000000000000000000));
	assign quotient_raw[3] = (~adder3_out[34] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder3_out[34:0] == 35'b00000000000000000000000000000000000));
	assign quotient_new[1] = quotient_raw[3] | quotient_raw[2];
	assign quotient_new[0] = quotient_raw[3] | (~quotient_raw[2] & quotient_raw[1]);
	assign twos_comp_b_sel = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign twos_comp_q_sel = ((~valid_ff & ~rem_ff) & (dividend_sign_ff ^ divisor_sign_ff)) & ~by_zero_case_ff;
	assign twos_comp_in[31:0] = ({32 {twos_comp_q_sel}} & q_ff[31:0]) | ({32 {twos_comp_b_sel}} & b_ff[31:0]);
	rvtwoscomp #(.WIDTH(32)) i_twos_comp(
		.din(twos_comp_in[31:0]),
		.dout(twos_comp_out[31:0])
	);
	assign valid_out = finish_ff & ~cancel;
	assign data_out[31:0] = (({32 {~rem_ff & ~twos_comp_q_sel}} & q_ff[31:0]) | ({32 {rem_ff}} & r_ff[31:0])) | ({32 {twos_comp_q_sel}} & twos_comp_out[31:0]);
	assign smallnum_case = ((((((a_ff[31:4] == 28'b0000000000000000000000000000) & (b_ff[31:4] == 28'b0000000000000000000000000000)) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel) | (((((a_ff[31:0] == 32'b00000000000000000000000000000000) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel);
	assign smallnum[3] = ((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1];
	assign smallnum[2] = ((((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[2]);
	assign smallnum[1] = ((((((((((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[1]) & ~b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]);
	assign smallnum[0] = ((((((((((((((((((((((((((((a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1]) | (((((a_ff[3] & ~a_ff[2]) & a_ff[0]) & ~b_ff[3]) & b_ff[1]) & b_ff[0])) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0])) | (((a_ff[0] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | ((((((~a_ff[3] & a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[0])) | (((a_ff[3] & ~b_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | ((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & b_ff[2]) & b_ff[1])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | ((((~a_ff[3] & a_ff[2]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[0])) | ((((~a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[3] & a_ff[1]) & ~b_ff[2]) & ~b_ff[0])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & b_ff[2])) | (((a_ff[3] & a_ff[2]) & b_ff[3]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[1]) & b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[0]) & ~b_ff[2]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[0]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & ~a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[1])) | (((a_ff[3] & a_ff[1]) & a_ff[0]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & b_ff[3]);
	assign shortq_dividend[32:0] = {dividend_sign_ff, a_ff[31:0]};
	wire [5:0] dw_a_enc;
	wire [5:0] dw_b_enc;
	wire [6:0] dw_shortq_raw;
	eb1_exu_div_cls i_a_cls(
		.operand(shortq_dividend[32:0]),
		.cls(dw_a_enc[4:0])
	);
	eb1_exu_div_cls i_b_cls(
		.operand(b_ff[32:0]),
		.cls(dw_b_enc[4:0])
	);
	assign dw_a_enc[5] = 1'b0;
	assign dw_b_enc[5] = 1'b0;
	assign dw_shortq_raw[6:0] = ({1'b0, dw_b_enc[5:0]} - {1'b0, dw_a_enc[5:0]}) + 7'd1;
	assign shortq[5:0] = (dw_shortq_raw[6] ? 6'd0 : dw_shortq_raw[5:0]);
	assign shortq_enable = ((valid_ff & ~shortq[5]) & ~(shortq[4:1] == 4'b1111)) & ~cancel;
	assign shortq_shift[4:0] = (~shortq_enable ? 5'd0 : 5'b11111 - shortq[4:0]);
endmodule
module eb1_exu_div_new_3bit_fullshortq (
	clk,
	rst_l,
	scan_mode,
	cancel,
	valid_in,
	signed_in,
	rem_in,
	dividend_in,
	divisor_in,
	valid_out,
	data_out
);
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire cancel;
	input wire valid_in;
	input wire signed_in;
	input wire rem_in;
	input wire [31:0] dividend_in;
	input wire [31:0] divisor_in;
	output wire valid_out;
	output wire [31:0] data_out;
	wire valid_ff_in;
	wire valid_ff;
	wire finish_raw;
	wire finish;
	wire finish_ff;
	wire running_state;
	wire misc_enable;
	wire [2:0] control_in;
	wire [2:0] control_ff;
	wire dividend_sign_ff;
	wire divisor_sign_ff;
	wire rem_ff;
	wire count_enable;
	wire [6:0] count_in;
	wire [6:0] count_ff;
	wire smallnum_case;
	wire [3:0] smallnum;
	wire a_enable;
	wire a_shift;
	wire [32:0] a_in;
	wire [32:0] a_ff;
	wire b_enable;
	wire b_twos_comp;
	wire [32:0] b_in;
	wire [36:0] b_ff;
	wire [31:0] q_in;
	wire [31:0] q_ff;
	wire rq_enable;
	wire r_sign_sel;
	wire r_restore_sel;
	wire r_adder1_sel;
	wire r_adder2_sel;
	wire r_adder3_sel;
	wire r_adder4_sel;
	wire r_adder5_sel;
	wire r_adder6_sel;
	wire r_adder7_sel;
	wire [32:0] r_in;
	wire [32:0] r_ff;
	wire twos_comp_q_sel;
	wire twos_comp_b_sel;
	wire [31:0] twos_comp_in;
	wire [31:0] twos_comp_out;
	wire [7:1] quotient_raw;
	wire [2:0] quotient_new;
	wire [33:0] adder1_out;
	wire [34:0] adder2_out;
	wire [35:0] adder3_out;
	wire [36:0] adder4_out;
	wire [36:0] adder5_out;
	wire [36:0] adder6_out;
	wire [36:0] adder7_out;
	wire [65:0] ar_shifted;
	wire [5:0] shortq;
	wire [4:0] shortq_shift;
	wire [4:0] shortq_decode;
	wire [4:0] shortq_shift_ff;
	wire shortq_enable;
	wire shortq_enable_ff;
	wire [32:0] shortq_dividend;
	wire by_zero_case;
	wire by_zero_case_ff;
	rvdffe #(.WIDTH(19)) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(misc_enable),
		.din({valid_ff_in, control_in[2:0], by_zero_case, shortq_enable, shortq_shift[4:0], finish, count_in[6:0]}),
		.dout({valid_ff, control_ff[2:0], by_zero_case_ff, shortq_enable_ff, shortq_shift_ff[4:0], finish_ff, count_ff[6:0]})
	);
	rvdffe #(.WIDTH(33)) i_a_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(a_enable),
		.din(a_in[32:0]),
		.dout(a_ff[32:0])
	);
	rvdffe #(.WIDTH(33)) i_b_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(b_enable),
		.din(b_in[32:0]),
		.dout(b_ff[32:0])
	);
	rvdffe #(.WIDTH(33)) i_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(r_in[32:0]),
		.dout(r_ff[32:0])
	);
	rvdffe #(.WIDTH(32)) i_q_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(q_in[31:0]),
		.dout(q_ff[31:0])
	);
	assign valid_ff_in = valid_in & ~cancel;
	assign control_in[2] = (~valid_in & control_ff[2]) | ((valid_in & signed_in) & dividend_in[31]);
	assign control_in[1] = (~valid_in & control_ff[1]) | ((valid_in & signed_in) & divisor_in[31]);
	assign control_in[0] = (~valid_in & control_ff[0]) | (valid_in & rem_in);
	assign dividend_sign_ff = control_ff[2];
	assign divisor_sign_ff = control_ff[1];
	assign rem_ff = control_ff[0];
	assign by_zero_case = valid_ff & (b_ff[31:0] == 32'b00000000000000000000000000000000);
	assign misc_enable = (((valid_in | valid_ff) | cancel) | running_state) | finish_ff;
	assign running_state = |count_ff[6:0] | shortq_enable_ff;
	assign finish_raw = (smallnum_case | by_zero_case) | (count_ff[6:0] == 7'd33);
	assign finish = finish_raw & ~cancel;
	assign count_enable = ((((valid_ff | running_state) & ~finish) & ~finish_ff) & ~cancel) & ~shortq_enable;
	assign count_in[6:0] = {7 {count_enable}} & ((count_ff[6:0] + 7'b0000011) + {2'b00, shortq_shift_ff[4:0]});
	assign a_enable = valid_in | running_state;
	assign a_shift = running_state & ~shortq_enable_ff;
	assign ar_shifted[65:0] = {{33 {dividend_sign_ff}}, a_ff[32:0]} << {shortq_shift_ff[4:0]};
	assign a_in[32:0] = (({33 {~a_shift & ~shortq_enable_ff}} & {signed_in & dividend_in[31], dividend_in[31:0]}) | ({33 {a_shift}} & {a_ff[29:0], 3'b000})) | ({33 {shortq_enable_ff}} & ar_shifted[32:0]);
	assign b_enable = valid_in | b_twos_comp;
	assign b_twos_comp = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign b_in[32:0] = ({33 {~b_twos_comp}} & {signed_in & divisor_in[31], divisor_in[31:0]}) | ({33 {b_twos_comp}} & {~divisor_sign_ff, twos_comp_out[31:0]});
	assign rq_enable = (valid_in | valid_ff) | running_state;
	assign r_sign_sel = (valid_ff & dividend_sign_ff) & ~by_zero_case;
	assign r_restore_sel = (running_state & (quotient_new[2:0] == 3'b000)) & ~shortq_enable_ff;
	assign r_adder1_sel = (running_state & (quotient_new[2:0] == 3'b001)) & ~shortq_enable_ff;
	assign r_adder2_sel = (running_state & (quotient_new[2:0] == 3'b010)) & ~shortq_enable_ff;
	assign r_adder3_sel = (running_state & (quotient_new[2:0] == 3'b011)) & ~shortq_enable_ff;
	assign r_adder4_sel = (running_state & (quotient_new[2:0] == 3'b100)) & ~shortq_enable_ff;
	assign r_adder5_sel = (running_state & (quotient_new[2:0] == 3'b101)) & ~shortq_enable_ff;
	assign r_adder6_sel = (running_state & (quotient_new[2:0] == 3'b110)) & ~shortq_enable_ff;
	assign r_adder7_sel = (running_state & (quotient_new[2:0] == 3'b111)) & ~shortq_enable_ff;
	assign r_in[32:0] = (((((((((({33 {r_sign_sel}} & {33 {1'b1}}) | ({33 {r_restore_sel}} & {r_ff[29:0], a_ff[32:30]})) | ({33 {r_adder1_sel}} & adder1_out[32:0])) | ({33 {r_adder2_sel}} & adder2_out[32:0])) | ({33 {r_adder3_sel}} & adder3_out[32:0])) | ({33 {r_adder4_sel}} & adder4_out[32:0])) | ({33 {r_adder5_sel}} & adder5_out[32:0])) | ({33 {r_adder6_sel}} & adder6_out[32:0])) | ({33 {r_adder7_sel}} & adder7_out[32:0])) | ({33 {shortq_enable_ff}} & ar_shifted[65:33])) | ({33 {by_zero_case}} & {1'b0, a_ff[31:0]});
	assign q_in[31:0] = (({32 {~valid_ff}} & {q_ff[28:0], quotient_new[2:0]}) | ({32 {smallnum_case}} & {28'b0000000000000000000000000000, smallnum[3:0]})) | ({32 {by_zero_case}} & {32 {1'b1}});
	assign b_ff[36:33] = {b_ff[32], b_ff[32], b_ff[32], b_ff[32]};
	assign adder1_out[33:0] = {r_ff[30:0], a_ff[32:30]} + b_ff[33:0];
	assign adder2_out[34:0] = {r_ff[31:0], a_ff[32:30]} + {b_ff[33:0], 1'b0};
	assign adder3_out[35:0] = ({r_ff[32:0], a_ff[32:30]} + {b_ff[34:0], 1'b0}) + b_ff[35:0];
	assign adder4_out[36:0] = {r_ff[32], r_ff[32:0], a_ff[32:30]} + {b_ff[34:0], 2'b00};
	assign adder5_out[36:0] = ({r_ff[32], r_ff[32:0], a_ff[32:30]} + {b_ff[34:0], 2'b00}) + b_ff[36:0];
	assign adder6_out[36:0] = ({r_ff[32], r_ff[32:0], a_ff[32:30]} + {b_ff[34:0], 2'b00}) + {b_ff[35:0], 1'b0};
	assign adder7_out[36:0] = (({r_ff[32], r_ff[32:0], a_ff[32:30]} + {b_ff[34:0], 2'b00}) + {b_ff[35:0], 1'b0}) + b_ff[36:0];
	assign quotient_raw[1] = (~adder1_out[33] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder1_out[33:0] == 34'b0000000000000000000000000000000000));
	assign quotient_raw[2] = (~adder2_out[34] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder2_out[34:0] == 35'b00000000000000000000000000000000000));
	assign quotient_raw[3] = (~adder3_out[35] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder3_out[35:0] == 36'b000000000000000000000000000000000000));
	assign quotient_raw[4] = (~adder4_out[36] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder4_out[36:0] == 37'b0000000000000000000000000000000000000));
	assign quotient_raw[5] = (~adder5_out[36] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder5_out[36:0] == 37'b0000000000000000000000000000000000000));
	assign quotient_raw[6] = (~adder6_out[36] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder6_out[36:0] == 37'b0000000000000000000000000000000000000));
	assign quotient_raw[7] = (~adder7_out[36] ^ dividend_sign_ff) | ((a_ff[29:0] == 30'b000000000000000000000000000000) & (adder7_out[36:0] == 37'b0000000000000000000000000000000000000));
	assign quotient_new[2] = ((quotient_raw[7] | quotient_raw[6]) | quotient_raw[5]) | quotient_raw[4];
	assign quotient_new[1] = ((quotient_raw[7] | quotient_raw[6]) | (~quotient_raw[4] & quotient_raw[3])) | (~quotient_raw[3] & quotient_raw[2]);
	assign quotient_new[0] = ((quotient_raw[7] | (~quotient_raw[6] & quotient_raw[5])) | (~quotient_raw[4] & quotient_raw[3])) | (~quotient_raw[2] & quotient_raw[1]);
	assign twos_comp_b_sel = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign twos_comp_q_sel = ((~valid_ff & ~rem_ff) & (dividend_sign_ff ^ divisor_sign_ff)) & ~by_zero_case_ff;
	assign twos_comp_in[31:0] = ({32 {twos_comp_q_sel}} & q_ff[31:0]) | ({32 {twos_comp_b_sel}} & b_ff[31:0]);
	rvtwoscomp #(.WIDTH(32)) i_twos_comp(
		.din(twos_comp_in[31:0]),
		.dout(twos_comp_out[31:0])
	);
	assign valid_out = finish_ff & ~cancel;
	assign data_out[31:0] = (({32 {~rem_ff & ~twos_comp_q_sel}} & q_ff[31:0]) | ({32 {rem_ff}} & r_ff[31:0])) | ({32 {twos_comp_q_sel}} & twos_comp_out[31:0]);
	assign smallnum_case = ((((((a_ff[31:4] == 28'b0000000000000000000000000000) & (b_ff[31:4] == 28'b0000000000000000000000000000)) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel) | (((((a_ff[31:0] == 32'b00000000000000000000000000000000) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel);
	assign smallnum[3] = ((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1];
	assign smallnum[2] = ((((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[2]);
	assign smallnum[1] = ((((((((((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[1]) & ~b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]);
	assign smallnum[0] = ((((((((((((((((((((((((((((a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1]) | (((((a_ff[3] & ~a_ff[2]) & a_ff[0]) & ~b_ff[3]) & b_ff[1]) & b_ff[0])) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0])) | (((a_ff[0] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | ((((((~a_ff[3] & a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[0])) | (((a_ff[3] & ~b_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | ((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & b_ff[2]) & b_ff[1])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | ((((~a_ff[3] & a_ff[2]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[0])) | ((((~a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[3] & a_ff[1]) & ~b_ff[2]) & ~b_ff[0])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & b_ff[2])) | (((a_ff[3] & a_ff[2]) & b_ff[3]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[1]) & b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[0]) & ~b_ff[2]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[0]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & ~a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[1])) | (((a_ff[3] & a_ff[1]) & a_ff[0]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & b_ff[3]);
	assign shortq_dividend[32:0] = {dividend_sign_ff, a_ff[31:0]};
	wire [5:0] dw_a_enc;
	wire [5:0] dw_b_enc;
	wire [6:0] dw_shortq_raw;
	eb1_exu_div_cls i_a_cls(
		.operand(shortq_dividend[32:0]),
		.cls(dw_a_enc[4:0])
	);
	eb1_exu_div_cls i_b_cls(
		.operand(b_ff[32:0]),
		.cls(dw_b_enc[4:0])
	);
	assign dw_a_enc[5] = 1'b0;
	assign dw_b_enc[5] = 1'b0;
	assign dw_shortq_raw[6:0] = ({1'b0, dw_b_enc[5:0]} - {1'b0, dw_a_enc[5:0]}) + 7'd1;
	assign shortq[5:0] = (dw_shortq_raw[6] ? 6'd0 : dw_shortq_raw[5:0]);
	assign shortq_enable = ((valid_ff & ~shortq[5]) & ~(shortq[4:2] == 3'b111)) & ~cancel;
	assign shortq_decode[4:0] = ((((((((((((((((((((((((((((((({5 {shortq[4:0] == 5'd31}} & 5'd0) | ({5 {shortq[4:0] == 5'd30}} & 5'd0)) | ({5 {shortq[4:0] == 5'd29}} & 5'd0)) | ({5 {shortq[4:0] == 5'd28}} & 5'd0)) | ({5 {shortq[4:0] == 5'd27}} & 5'd3)) | ({5 {shortq[4:0] == 5'd26}} & 5'd6)) | ({5 {shortq[4:0] == 5'd25}} & 5'd6)) | ({5 {shortq[4:0] == 5'd24}} & 5'd6)) | ({5 {shortq[4:0] == 5'd23}} & 5'd9)) | ({5 {shortq[4:0] == 5'd22}} & 5'd9)) | ({5 {shortq[4:0] == 5'd21}} & 5'd9)) | ({5 {shortq[4:0] == 5'd20}} & 5'd12)) | ({5 {shortq[4:0] == 5'd19}} & 5'd12)) | ({5 {shortq[4:0] == 5'd18}} & 5'd12)) | ({5 {shortq[4:0] == 5'd17}} & 5'd15)) | ({5 {shortq[4:0] == 5'd16}} & 5'd15)) | ({5 {shortq[4:0] == 5'd15}} & 5'd15)) | ({5 {shortq[4:0] == 5'd14}} & 5'd18)) | ({5 {shortq[4:0] == 5'd13}} & 5'd18)) | ({5 {shortq[4:0] == 5'd12}} & 5'd18)) | ({5 {shortq[4:0] == 5'd11}} & 5'd21)) | ({5 {shortq[4:0] == 5'd10}} & 5'd21)) | ({5 {shortq[4:0] == 5'd9}} & 5'd21)) | ({5 {shortq[4:0] == 5'd8}} & 5'd24)) | ({5 {shortq[4:0] == 5'd7}} & 5'd24)) | ({5 {shortq[4:0] == 5'd6}} & 5'd24)) | ({5 {shortq[4:0] == 5'd5}} & 5'd27)) | ({5 {shortq[4:0] == 5'd4}} & 5'd27)) | ({5 {shortq[4:0] == 5'd3}} & 5'd27)) | ({5 {shortq[4:0] == 5'd2}} & 5'd27)) | ({5 {shortq[4:0] == 5'd1}} & 5'd27)) | ({5 {shortq[4:0] == 5'd0}} & 5'd27);
	assign shortq_shift[4:0] = (~shortq_enable ? 5'd0 : shortq_decode[4:0]);
endmodule
module eb1_exu_div_new_4bit_fullshortq (
	clk,
	rst_l,
	scan_mode,
	cancel,
	valid_in,
	signed_in,
	rem_in,
	dividend_in,
	divisor_in,
	valid_out,
	data_out
);
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire cancel;
	input wire valid_in;
	input wire signed_in;
	input wire rem_in;
	input wire [31:0] dividend_in;
	input wire [31:0] divisor_in;
	output wire valid_out;
	output wire [31:0] data_out;
	wire valid_ff_in;
	wire valid_ff;
	wire finish_raw;
	wire finish;
	wire finish_ff;
	wire running_state;
	wire misc_enable;
	wire [2:0] control_in;
	wire [2:0] control_ff;
	wire dividend_sign_ff;
	wire divisor_sign_ff;
	wire rem_ff;
	wire count_enable;
	wire [6:0] count_in;
	wire [6:0] count_ff;
	wire smallnum_case;
	wire [3:0] smallnum;
	wire a_enable;
	wire a_shift;
	wire [31:0] a_in;
	wire [31:0] a_ff;
	wire b_enable;
	wire b_twos_comp;
	wire [32:0] b_in;
	wire [37:0] b_ff;
	wire [31:0] q_in;
	wire [31:0] q_ff;
	wire rq_enable;
	wire r_sign_sel;
	wire r_restore_sel;
	wire r_adder01_sel;
	wire r_adder02_sel;
	wire r_adder03_sel;
	wire r_adder04_sel;
	wire r_adder05_sel;
	wire r_adder06_sel;
	wire r_adder07_sel;
	wire r_adder08_sel;
	wire r_adder09_sel;
	wire r_adder10_sel;
	wire r_adder11_sel;
	wire r_adder12_sel;
	wire r_adder13_sel;
	wire r_adder14_sel;
	wire r_adder15_sel;
	wire [32:0] r_in;
	wire [32:0] r_ff;
	wire twos_comp_q_sel;
	wire twos_comp_b_sel;
	wire [31:0] twos_comp_in;
	wire [31:0] twos_comp_out;
	wire [15:1] quotient_raw;
	wire [3:0] quotient_new;
	wire [34:0] adder01_out;
	wire [35:0] adder02_out;
	wire [36:0] adder03_out;
	wire [37:0] adder04_out;
	wire [37:0] adder05_out;
	wire [37:0] adder06_out;
	wire [37:0] adder07_out;
	wire [37:0] adder08_out;
	wire [37:0] adder09_out;
	wire [37:0] adder10_out;
	wire [37:0] adder11_out;
	wire [37:0] adder12_out;
	wire [37:0] adder13_out;
	wire [37:0] adder14_out;
	wire [37:0] adder15_out;
	wire [64:0] ar_shifted;
	wire [5:0] shortq;
	wire [4:0] shortq_shift;
	wire [4:0] shortq_decode;
	wire [4:0] shortq_shift_ff;
	wire shortq_enable;
	wire shortq_enable_ff;
	wire [32:0] shortq_dividend;
	wire by_zero_case;
	wire by_zero_case_ff;
	rvdffe #(.WIDTH(19)) i_misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(misc_enable),
		.din({valid_ff_in, control_in[2:0], by_zero_case, shortq_enable, shortq_shift[4:0], finish, count_in[6:0]}),
		.dout({valid_ff, control_ff[2:0], by_zero_case_ff, shortq_enable_ff, shortq_shift_ff[4:0], finish_ff, count_ff[6:0]})
	);
	rvdffe #(.WIDTH(32)) i_a_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(a_enable),
		.din(a_in[31:0]),
		.dout(a_ff[31:0])
	);
	rvdffe #(.WIDTH(33)) i_b_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(b_enable),
		.din(b_in[32:0]),
		.dout(b_ff[32:0])
	);
	rvdffe #(.WIDTH(33)) i_r_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(r_in[32:0]),
		.dout(r_ff[32:0])
	);
	rvdffe #(.WIDTH(32)) i_q_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(rq_enable),
		.din(q_in[31:0]),
		.dout(q_ff[31:0])
	);
	assign valid_ff_in = valid_in & ~cancel;
	assign control_in[2] = (~valid_in & control_ff[2]) | ((valid_in & signed_in) & dividend_in[31]);
	assign control_in[1] = (~valid_in & control_ff[1]) | ((valid_in & signed_in) & divisor_in[31]);
	assign control_in[0] = (~valid_in & control_ff[0]) | (valid_in & rem_in);
	assign dividend_sign_ff = control_ff[2];
	assign divisor_sign_ff = control_ff[1];
	assign rem_ff = control_ff[0];
	assign by_zero_case = valid_ff & (b_ff[31:0] == 32'b00000000000000000000000000000000);
	assign misc_enable = (((valid_in | valid_ff) | cancel) | running_state) | finish_ff;
	assign running_state = |count_ff[6:0] | shortq_enable_ff;
	assign finish_raw = (smallnum_case | by_zero_case) | (count_ff[6:0] == 7'd32);
	assign finish = finish_raw & ~cancel;
	assign count_enable = ((((valid_ff | running_state) & ~finish) & ~finish_ff) & ~cancel) & ~shortq_enable;
	assign count_in[6:0] = {7 {count_enable}} & ((count_ff[6:0] + 7'd4) + {2'b00, shortq_shift_ff[4:0]});
	assign a_enable = valid_in | running_state;
	assign a_shift = running_state & ~shortq_enable_ff;
	assign ar_shifted[64:0] = {{33 {dividend_sign_ff}}, a_ff[31:0]} << {shortq_shift_ff[4:0]};
	assign a_in[31:0] = (({32 {~a_shift & ~shortq_enable_ff}} & dividend_in[31:0]) | ({32 {a_shift}} & {a_ff[27:0], 4'b0000})) | ({32 {shortq_enable_ff}} & ar_shifted[31:0]);
	assign b_enable = valid_in | b_twos_comp;
	assign b_twos_comp = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign b_in[32:0] = ({33 {~b_twos_comp}} & {signed_in & divisor_in[31], divisor_in[31:0]}) | ({33 {b_twos_comp}} & {~divisor_sign_ff, twos_comp_out[31:0]});
	assign rq_enable = (valid_in | valid_ff) | running_state;
	assign r_sign_sel = (valid_ff & dividend_sign_ff) & ~by_zero_case;
	assign r_restore_sel = (running_state & (quotient_new[3:0] == 4'd0)) & ~shortq_enable_ff;
	assign r_adder01_sel = (running_state & (quotient_new[3:0] == 4'd1)) & ~shortq_enable_ff;
	assign r_adder02_sel = (running_state & (quotient_new[3:0] == 4'd2)) & ~shortq_enable_ff;
	assign r_adder03_sel = (running_state & (quotient_new[3:0] == 4'd3)) & ~shortq_enable_ff;
	assign r_adder04_sel = (running_state & (quotient_new[3:0] == 4'd4)) & ~shortq_enable_ff;
	assign r_adder05_sel = (running_state & (quotient_new[3:0] == 4'd5)) & ~shortq_enable_ff;
	assign r_adder06_sel = (running_state & (quotient_new[3:0] == 4'd6)) & ~shortq_enable_ff;
	assign r_adder07_sel = (running_state & (quotient_new[3:0] == 4'd7)) & ~shortq_enable_ff;
	assign r_adder08_sel = (running_state & (quotient_new[3:0] == 4'd8)) & ~shortq_enable_ff;
	assign r_adder09_sel = (running_state & (quotient_new[3:0] == 4'd9)) & ~shortq_enable_ff;
	assign r_adder10_sel = (running_state & (quotient_new[3:0] == 4'd10)) & ~shortq_enable_ff;
	assign r_adder11_sel = (running_state & (quotient_new[3:0] == 4'd11)) & ~shortq_enable_ff;
	assign r_adder12_sel = (running_state & (quotient_new[3:0] == 4'd12)) & ~shortq_enable_ff;
	assign r_adder13_sel = (running_state & (quotient_new[3:0] == 4'd13)) & ~shortq_enable_ff;
	assign r_adder14_sel = (running_state & (quotient_new[3:0] == 4'd14)) & ~shortq_enable_ff;
	assign r_adder15_sel = (running_state & (quotient_new[3:0] == 4'd15)) & ~shortq_enable_ff;
	assign r_in[32:0] = (((((((((((((((((({33 {r_sign_sel}} & {33 {1'b1}}) | ({33 {r_restore_sel}} & {r_ff[28:0], a_ff[31:28]})) | ({33 {r_adder01_sel}} & adder01_out[32:0])) | ({33 {r_adder02_sel}} & adder02_out[32:0])) | ({33 {r_adder03_sel}} & adder03_out[32:0])) | ({33 {r_adder04_sel}} & adder04_out[32:0])) | ({33 {r_adder05_sel}} & adder05_out[32:0])) | ({33 {r_adder06_sel}} & adder06_out[32:0])) | ({33 {r_adder07_sel}} & adder07_out[32:0])) | ({33 {r_adder08_sel}} & adder08_out[32:0])) | ({33 {r_adder09_sel}} & adder09_out[32:0])) | ({33 {r_adder10_sel}} & adder10_out[32:0])) | ({33 {r_adder11_sel}} & adder11_out[32:0])) | ({33 {r_adder12_sel}} & adder12_out[32:0])) | ({33 {r_adder13_sel}} & adder13_out[32:0])) | ({33 {r_adder14_sel}} & adder14_out[32:0])) | ({33 {r_adder15_sel}} & adder15_out[32:0])) | ({33 {shortq_enable_ff}} & ar_shifted[64:32])) | ({33 {by_zero_case}} & {1'b0, a_ff[31:0]});
	assign q_in[31:0] = (({32 {~valid_ff}} & {q_ff[27:0], quotient_new[3:0]}) | ({32 {smallnum_case}} & {28'b0000000000000000000000000000, smallnum[3:0]})) | ({32 {by_zero_case}} & {32 {1'b1}});
	assign b_ff[37:33] = {b_ff[32], b_ff[32], b_ff[32], b_ff[32], b_ff[32]};
	assign adder01_out[34:0] = {r_ff[30:0], a_ff[31:28]} + b_ff[34:0];
	assign adder02_out[35:0] = {r_ff[31:0], a_ff[31:28]} + {b_ff[34:0], 1'b0};
	assign adder03_out[36:0] = ({r_ff[32:0], a_ff[31:28]} + {b_ff[35:0], 1'b0}) + b_ff[36:0];
	assign adder04_out[37:0] = {r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[35:0], 2'b00};
	assign adder05_out[37:0] = ({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[35:0], 2'b00}) + b_ff[37:0];
	assign adder06_out[37:0] = ({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[35:0], 2'b00}) + {b_ff[36:0], 1'b0};
	assign adder07_out[37:0] = (({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[35:0], 2'b00}) + {b_ff[36:0], 1'b0}) + b_ff[37:0];
	assign adder08_out[37:0] = {r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000};
	assign adder09_out[37:0] = ({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + b_ff[37:0];
	assign adder10_out[37:0] = ({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[36:0], 1'b0};
	assign adder11_out[37:0] = (({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[36:0], 1'b0}) + b_ff[37:0];
	assign adder12_out[37:0] = ({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[35:0], 2'b00};
	assign adder13_out[37:0] = (({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[35:0], 2'b00}) + b_ff[37:0];
	assign adder14_out[37:0] = (({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[35:0], 2'b00}) + {b_ff[36:0], 1'b0};
	assign adder15_out[37:0] = ((({r_ff[32], r_ff[32:0], a_ff[31:28]} + {b_ff[34:0], 3'b000}) + {b_ff[35:0], 2'b00}) + {b_ff[36:0], 1'b0}) + b_ff[37:0];
	assign quotient_raw[1] = (~adder01_out[34] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder01_out[34:0] == 35'b00000000000000000000000000000000000));
	assign quotient_raw[2] = (~adder02_out[35] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder02_out[35:0] == 36'b000000000000000000000000000000000000));
	assign quotient_raw[3] = (~adder03_out[36] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder03_out[36:0] == 37'b0000000000000000000000000000000000000));
	assign quotient_raw[4] = (~adder04_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder04_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[5] = (~adder05_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder05_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[6] = (~adder06_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder06_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[7] = (~adder07_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder07_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[8] = (~adder08_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder08_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[9] = (~adder09_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder09_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[10] = (~adder10_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder10_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[11] = (~adder11_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder11_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[12] = (~adder12_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder12_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[13] = (~adder13_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder13_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[14] = (~adder14_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder14_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_raw[15] = (~adder15_out[37] ^ dividend_sign_ff) | ((a_ff[27:0] == 28'b0000000000000000000000000000) & (adder15_out[37:0] == 38'b00000000000000000000000000000000000000));
	assign quotient_new[0] = (((((((quotient_raw[15:1] == 15'b000000000000001) | (quotient_raw[15:3] == 13'b0000000000001)) | (quotient_raw[15:5] == 11'b00000000001)) | (quotient_raw[15:7] == 9'b000000001)) | (quotient_raw[15:9] == 7'b0000001)) | (quotient_raw[15:11] == 5'b00001)) | (quotient_raw[15:13] == 3'b001)) | (quotient_raw[15] == 1'b1);
	assign quotient_new[1] = (((((((quotient_raw[15:2] == 14'b00000000000001) | (quotient_raw[15:3] == 13'b0000000000001)) | (quotient_raw[15:6] == 10'b0000000001)) | (quotient_raw[15:7] == 9'b000000001)) | (quotient_raw[15:10] == 6'b000001)) | (quotient_raw[15:11] == 5'b00001)) | (quotient_raw[15:14] == 2'b01)) | (quotient_raw[15] == 1'b1);
	assign quotient_new[2] = (((((((quotient_raw[15:4] == 12'b000000000001) | (quotient_raw[15:5] == 11'b00000000001)) | (quotient_raw[15:6] == 10'b0000000001)) | (quotient_raw[15:7] == 9'b000000001)) | (quotient_raw[15:12] == 4'b0001)) | (quotient_raw[15:13] == 3'b001)) | (quotient_raw[15:14] == 2'b01)) | (quotient_raw[15] == 1'b1);
	assign quotient_new[3] = (((((((quotient_raw[15:8] == 8'b00000001) | (quotient_raw[15:9] == 7'b0000001)) | (quotient_raw[15:10] == 6'b000001)) | (quotient_raw[15:11] == 5'b00001)) | (quotient_raw[15:12] == 4'b0001)) | (quotient_raw[15:13] == 3'b001)) | (quotient_raw[15:14] == 2'b01)) | (quotient_raw[15] == 1'b1);
	assign twos_comp_b_sel = valid_ff & ~(dividend_sign_ff ^ divisor_sign_ff);
	assign twos_comp_q_sel = ((~valid_ff & ~rem_ff) & (dividend_sign_ff ^ divisor_sign_ff)) & ~by_zero_case_ff;
	assign twos_comp_in[31:0] = ({32 {twos_comp_q_sel}} & q_ff[31:0]) | ({32 {twos_comp_b_sel}} & b_ff[31:0]);
	rvtwoscomp #(.WIDTH(32)) i_twos_comp(
		.din(twos_comp_in[31:0]),
		.dout(twos_comp_out[31:0])
	);
	assign valid_out = finish_ff & ~cancel;
	assign data_out[31:0] = (({32 {~rem_ff & ~twos_comp_q_sel}} & q_ff[31:0]) | ({32 {rem_ff}} & r_ff[31:0])) | ({32 {twos_comp_q_sel}} & twos_comp_out[31:0]);
	assign smallnum_case = ((((((a_ff[31:4] == 28'b0000000000000000000000000000) & (b_ff[31:4] == 28'b0000000000000000000000000000)) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel) | (((((a_ff[31:0] == 32'b00000000000000000000000000000000) & ~by_zero_case) & ~rem_ff) & valid_ff) & ~cancel);
	assign smallnum[3] = ((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1];
	assign smallnum[2] = ((((a_ff[3] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[2]);
	assign smallnum[1] = ((((((((((a_ff[2] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0]) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[1]) & ~b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]);
	assign smallnum[0] = ((((((((((((((((((((((((((((a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1]) | (((((a_ff[3] & ~a_ff[2]) & a_ff[0]) & ~b_ff[3]) & b_ff[1]) & b_ff[0])) | (((a_ff[2] & ~b_ff[3]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[1] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[0])) | (((a_ff[0] & ~b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | ((((((~a_ff[3] & a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & ~b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & ~b_ff[0])) | (((a_ff[3] & ~b_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | ((((a_ff[3] & ~a_ff[2]) & ~b_ff[3]) & b_ff[2]) & b_ff[1])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[2]) & ~b_ff[1])) | ((((~a_ff[3] & a_ff[2]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[2]) & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[0])) | ((((~a_ff[2] & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & ~b_ff[2])) | (((a_ff[3] & a_ff[2]) & ~b_ff[1]) & ~b_ff[0])) | (((a_ff[3] & a_ff[1]) & ~b_ff[2]) & ~b_ff[0])) | (((((~a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & ~b_ff[3]) & b_ff[2])) | (((a_ff[3] & a_ff[2]) & b_ff[3]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[1]) & b_ff[3]) & ~b_ff[2]) & ~b_ff[1])) | (((a_ff[3] & a_ff[0]) & ~b_ff[2]) & ~b_ff[1])) | (((((a_ff[3] & ~a_ff[1]) & ~b_ff[3]) & b_ff[2]) & b_ff[1]) & b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[0])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & a_ff[2]) & a_ff[0]) & b_ff[3]) & ~b_ff[1])) | ((((a_ff[3] & ~a_ff[2]) & a_ff[1]) & ~b_ff[3]) & b_ff[1])) | (((a_ff[3] & a_ff[1]) & a_ff[0]) & ~b_ff[2])) | ((((a_ff[3] & a_ff[2]) & a_ff[1]) & a_ff[0]) & b_ff[3]);
	assign shortq_dividend[32:0] = {dividend_sign_ff, a_ff[31:0]};
	wire [5:0] dw_a_enc;
	wire [5:0] dw_b_enc;
	wire [6:0] dw_shortq_raw;
	eb1_exu_div_cls i_a_cls(
		.operand(shortq_dividend[32:0]),
		.cls(dw_a_enc[4:0])
	);
	eb1_exu_div_cls i_b_cls(
		.operand(b_ff[32:0]),
		.cls(dw_b_enc[4:0])
	);
	assign dw_a_enc[5] = 1'b0;
	assign dw_b_enc[5] = 1'b0;
	assign dw_shortq_raw[6:0] = ({1'b0, dw_b_enc[5:0]} - {1'b0, dw_a_enc[5:0]}) + 7'd1;
	assign shortq[5:0] = (dw_shortq_raw[6] ? 6'd0 : dw_shortq_raw[5:0]);
	assign shortq_enable = ((valid_ff & ~shortq[5]) & ~(shortq[4:2] == 3'b111)) & ~cancel;
	assign shortq_decode[4:0] = ((((((((((((((((((((((((((((((({5 {shortq[4:0] == 5'd31}} & 5'd0) | ({5 {shortq[4:0] == 5'd30}} & 5'd0)) | ({5 {shortq[4:0] == 5'd29}} & 5'd0)) | ({5 {shortq[4:0] == 5'd28}} & 5'd0)) | ({5 {shortq[4:0] == 5'd27}} & 5'd4)) | ({5 {shortq[4:0] == 5'd26}} & 5'd4)) | ({5 {shortq[4:0] == 5'd25}} & 5'd4)) | ({5 {shortq[4:0] == 5'd24}} & 5'd4)) | ({5 {shortq[4:0] == 5'd23}} & 5'd8)) | ({5 {shortq[4:0] == 5'd22}} & 5'd8)) | ({5 {shortq[4:0] == 5'd21}} & 5'd8)) | ({5 {shortq[4:0] == 5'd20}} & 5'd8)) | ({5 {shortq[4:0] == 5'd19}} & 5'd12)) | ({5 {shortq[4:0] == 5'd18}} & 5'd12)) | ({5 {shortq[4:0] == 5'd17}} & 5'd12)) | ({5 {shortq[4:0] == 5'd16}} & 5'd12)) | ({5 {shortq[4:0] == 5'd15}} & 5'd16)) | ({5 {shortq[4:0] == 5'd14}} & 5'd16)) | ({5 {shortq[4:0] == 5'd13}} & 5'd16)) | ({5 {shortq[4:0] == 5'd12}} & 5'd16)) | ({5 {shortq[4:0] == 5'd11}} & 5'd20)) | ({5 {shortq[4:0] == 5'd10}} & 5'd20)) | ({5 {shortq[4:0] == 5'd9}} & 5'd20)) | ({5 {shortq[4:0] == 5'd8}} & 5'd20)) | ({5 {shortq[4:0] == 5'd7}} & 5'd24)) | ({5 {shortq[4:0] == 5'd6}} & 5'd24)) | ({5 {shortq[4:0] == 5'd5}} & 5'd24)) | ({5 {shortq[4:0] == 5'd4}} & 5'd24)) | ({5 {shortq[4:0] == 5'd3}} & 5'd28)) | ({5 {shortq[4:0] == 5'd2}} & 5'd28)) | ({5 {shortq[4:0] == 5'd1}} & 5'd28)) | ({5 {shortq[4:0] == 5'd0}} & 5'd28);
	assign shortq_shift[4:0] = (~shortq_enable ? 5'd0 : shortq_decode[4:0]);
endmodule
module eb1_exu_div_cls (
	operand,
	cls
);
	input wire [32:0] operand;
	output wire [4:0] cls;
	wire [4:0] cls_zeros;
	wire [4:0] cls_ones;
	assign cls_zeros[4:0] = (((((((((((((((((((((((((((((((({5 {operand[31] == 1'b1}} & 5'd0) | ({5 {operand[31:30] == 2'b01}} & 5'd1)) | ({5 {operand[31:29] == {{2 {1'b0}}, 1'b1}}} & 5'd2)) | ({5 {operand[31:28] == {{3 {1'b0}}, 1'b1}}} & 5'd3)) | ({5 {operand[31:27] == {{4 {1'b0}}, 1'b1}}} & 5'd4)) | ({5 {operand[31:26] == {{5 {1'b0}}, 1'b1}}} & 5'd5)) | ({5 {operand[31:25] == {{6 {1'b0}}, 1'b1}}} & 5'd6)) | ({5 {operand[31:24] == {{7 {1'b0}}, 1'b1}}} & 5'd7)) | ({5 {operand[31:23] == {{8 {1'b0}}, 1'b1}}} & 5'd8)) | ({5 {operand[31:22] == {{9 {1'b0}}, 1'b1}}} & 5'd9)) | ({5 {operand[31:21] == {{10 {1'b0}}, 1'b1}}} & 5'd10)) | ({5 {operand[31:20] == {{11 {1'b0}}, 1'b1}}} & 5'd11)) | ({5 {operand[31:19] == {{12 {1'b0}}, 1'b1}}} & 5'd12)) | ({5 {operand[31:18] == {{13 {1'b0}}, 1'b1}}} & 5'd13)) | ({5 {operand[31:17] == {{14 {1'b0}}, 1'b1}}} & 5'd14)) | ({5 {operand[31:16] == {{15 {1'b0}}, 1'b1}}} & 5'd15)) | ({5 {operand[31:15] == {{16 {1'b0}}, 1'b1}}} & 5'd16)) | ({5 {operand[31:14] == {{17 {1'b0}}, 1'b1}}} & 5'd17)) | ({5 {operand[31:13] == {{18 {1'b0}}, 1'b1}}} & 5'd18)) | ({5 {operand[31:12] == {{19 {1'b0}}, 1'b1}}} & 5'd19)) | ({5 {operand[31:11] == {{20 {1'b0}}, 1'b1}}} & 5'd20)) | ({5 {operand[31:10] == {{21 {1'b0}}, 1'b1}}} & 5'd21)) | ({5 {operand[31:9] == {{22 {1'b0}}, 1'b1}}} & 5'd22)) | ({5 {operand[31:8] == {{23 {1'b0}}, 1'b1}}} & 5'd23)) | ({5 {operand[31:7] == {{24 {1'b0}}, 1'b1}}} & 5'd24)) | ({5 {operand[31:6] == {{25 {1'b0}}, 1'b1}}} & 5'd25)) | ({5 {operand[31:5] == {{26 {1'b0}}, 1'b1}}} & 5'd26)) | ({5 {operand[31:4] == {{27 {1'b0}}, 1'b1}}} & 5'd27)) | ({5 {operand[31:3] == {{28 {1'b0}}, 1'b1}}} & 5'd28)) | ({5 {operand[31:2] == {{29 {1'b0}}, 1'b1}}} & 5'd29)) | ({5 {operand[31:1] == {{30 {1'b0}}, 1'b1}}} & 5'd30)) | ({5 {operand[31:0] == {{31 {1'b0}}, 1'b1}}} & 5'd31)) | ({5 {operand[31:0] == {32 {1'b0}}}} & 5'd0);
	assign cls_ones[4:0] = ((((((((((((((((((((((((((((((({5 {operand[31:30] == 2'b10}} & 5'd0) | ({5 {operand[31:29] == {{2 {1'b1}}, 1'b0}}} & 5'd1)) | ({5 {operand[31:28] == {{3 {1'b1}}, 1'b0}}} & 5'd2)) | ({5 {operand[31:27] == {{4 {1'b1}}, 1'b0}}} & 5'd3)) | ({5 {operand[31:26] == {{5 {1'b1}}, 1'b0}}} & 5'd4)) | ({5 {operand[31:25] == {{6 {1'b1}}, 1'b0}}} & 5'd5)) | ({5 {operand[31:24] == {{7 {1'b1}}, 1'b0}}} & 5'd6)) | ({5 {operand[31:23] == {{8 {1'b1}}, 1'b0}}} & 5'd7)) | ({5 {operand[31:22] == {{9 {1'b1}}, 1'b0}}} & 5'd8)) | ({5 {operand[31:21] == {{10 {1'b1}}, 1'b0}}} & 5'd9)) | ({5 {operand[31:20] == {{11 {1'b1}}, 1'b0}}} & 5'd10)) | ({5 {operand[31:19] == {{12 {1'b1}}, 1'b0}}} & 5'd11)) | ({5 {operand[31:18] == {{13 {1'b1}}, 1'b0}}} & 5'd12)) | ({5 {operand[31:17] == {{14 {1'b1}}, 1'b0}}} & 5'd13)) | ({5 {operand[31:16] == {{15 {1'b1}}, 1'b0}}} & 5'd14)) | ({5 {operand[31:15] == {{16 {1'b1}}, 1'b0}}} & 5'd15)) | ({5 {operand[31:14] == {{17 {1'b1}}, 1'b0}}} & 5'd16)) | ({5 {operand[31:13] == {{18 {1'b1}}, 1'b0}}} & 5'd17)) | ({5 {operand[31:12] == {{19 {1'b1}}, 1'b0}}} & 5'd18)) | ({5 {operand[31:11] == {{20 {1'b1}}, 1'b0}}} & 5'd19)) | ({5 {operand[31:10] == {{21 {1'b1}}, 1'b0}}} & 5'd20)) | ({5 {operand[31:9] == {{22 {1'b1}}, 1'b0}}} & 5'd21)) | ({5 {operand[31:8] == {{23 {1'b1}}, 1'b0}}} & 5'd22)) | ({5 {operand[31:7] == {{24 {1'b1}}, 1'b0}}} & 5'd23)) | ({5 {operand[31:6] == {{25 {1'b1}}, 1'b0}}} & 5'd24)) | ({5 {operand[31:5] == {{26 {1'b1}}, 1'b0}}} & 5'd25)) | ({5 {operand[31:4] == {{27 {1'b1}}, 1'b0}}} & 5'd26)) | ({5 {operand[31:3] == {{28 {1'b1}}, 1'b0}}} & 5'd27)) | ({5 {operand[31:2] == {{29 {1'b1}}, 1'b0}}} & 5'd28)) | ({5 {operand[31:1] == {{30 {1'b1}}, 1'b0}}} & 5'd29)) | ({5 {operand[31:0] == {{31 {1'b1}}, 1'b0}}} & 5'd30)) | ({5 {operand[31:0] == {32 {1'b1}}}} & 5'd31);
	assign cls[4:0] = (operand[32] ? cls_ones[4:0] : cls_zeros[4:0]);
endmodule
module eb1_exu_mul_ctl (
	clk,
	rst_l,
	scan_mode,
	mul_p,
	rs1_in,
	rs2_in,
	result_x
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire [19:0] mul_p;
	input wire [31:0] rs1_in;
	input wire [31:0] rs2_in;
	output wire [31:0] result_x;
	wire mul_x_enable;
	wire bit_x_enable;
	wire signed [32:0] rs1_ext_in;
	wire signed [32:0] rs2_ext_in;
	wire [65:0] prod_x;
	wire low_x;
	wire bitmanip_sel_d;
	wire bitmanip_sel_x;
	wire [31:0] bitmanip_d;
	wire [31:0] bitmanip_x;
	wire ap_bext;
	wire ap_bdep;
	wire ap_clmul;
	wire ap_clmulh;
	wire ap_clmulr;
	wire ap_grev;
	wire ap_gorc;
	wire ap_shfl;
	wire ap_unshfl;
	wire ap_crc32_b;
	wire ap_crc32_h;
	wire ap_crc32_w;
	wire ap_crc32c_b;
	wire ap_crc32c_h;
	wire ap_crc32c_w;
	wire ap_bfp;
	generate
		if (pt[2197-:5] == 1) begin
			assign ap_bext = mul_p[15];
			assign ap_bdep = mul_p[14];
		end
		else begin
			assign ap_bext = 1'b0;
			assign ap_bdep = 1'b0;
		end
	endgenerate
	generate
		if (pt[2202-:5] == 1) begin
			assign ap_clmul = mul_p[13];
			assign ap_clmulh = mul_p[12];
			assign ap_clmulr = mul_p[11];
		end
		else begin
			assign ap_clmul = 1'b0;
			assign ap_clmulh = 1'b0;
			assign ap_clmulr = 1'b0;
		end
	endgenerate
	generate
		if (pt[2187-:5] == 1) begin
			assign ap_grev = mul_p[10];
			assign ap_gorc = mul_p[9];
			assign ap_shfl = mul_p[8];
			assign ap_unshfl = mul_p[7];
		end
		else begin
			assign ap_grev = 1'b0;
			assign ap_gorc = 1'b0;
			assign ap_shfl = 1'b0;
			assign ap_unshfl = 1'b0;
		end
	endgenerate
	generate
		if (pt[2182-:5] == 1) begin
			assign ap_crc32_b = mul_p[6];
			assign ap_crc32_h = mul_p[5];
			assign ap_crc32_w = mul_p[4];
			assign ap_crc32c_b = mul_p[3];
			assign ap_crc32c_h = mul_p[2];
			assign ap_crc32c_w = mul_p[1];
		end
		else begin
			assign ap_crc32_b = 1'b0;
			assign ap_crc32_h = 1'b0;
			assign ap_crc32_w = 1'b0;
			assign ap_crc32c_b = 1'b0;
			assign ap_crc32c_h = 1'b0;
			assign ap_crc32c_w = 1'b0;
		end
	endgenerate
	generate
		if (pt[2192-:5] == 1) begin
			assign ap_bfp = mul_p[0];
		end
		else assign ap_bfp = 1'b0;
	endgenerate
	assign mul_x_enable = mul_p[19];
	assign bit_x_enable = mul_p[19];
	assign rs1_ext_in[32] = mul_p[18] & rs1_in[31];
	assign rs2_ext_in[32] = mul_p[17] & rs2_in[31];
	assign rs1_ext_in[31:0] = rs1_in[31:0];
	assign rs2_ext_in[31:0] = rs2_in[31:0];
	wire signed [32:0] rs1_x;
	wire signed [32:0] rs2_x;
	rvdffe #(.WIDTH(34)) i_a_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din({mul_p[16], rs1_ext_in[32:0]}),
		.dout({low_x, rs1_x[32:0]}),
		.en(mul_x_enable)
	);
	rvdffe #(.WIDTH(33)) i_b_x_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din(rs2_ext_in[32:0]),
		.dout(rs2_x[32:0]),
		.en(mul_x_enable)
	);
	assign prod_x[65:0] = rs1_x * rs2_x;
	reg [31:0] bext_d;
	reg bext_test_bit_d;
	integer bext_i;
	integer bext_j;
	always @(*) begin
		bext_j = 0;
		bext_test_bit_d = 1'b0;
		bext_d[31:0] = 32'b00000000000000000000000000000000;
		for (bext_i = 0; bext_i < 32; bext_i = bext_i + 1)
			begin
				bext_test_bit_d = rs2_in[bext_i];
				if (bext_test_bit_d) begin
					bext_d[bext_j] = rs1_in[bext_i];
					bext_j = bext_j + 1;
				end
			end
	end
	reg [31:0] bdep_d;
	reg bdep_test_bit_d;
	integer bdep_i;
	integer bdep_j;
	always @(*) begin
		bdep_j = 0;
		bdep_test_bit_d = 1'b0;
		bdep_d[31:0] = 32'b00000000000000000000000000000000;
		for (bdep_i = 0; bdep_i < 32; bdep_i = bdep_i + 1)
			begin
				bdep_test_bit_d = rs2_in[bdep_i];
				if (bdep_test_bit_d) begin
					bdep_d[bdep_i] = rs1_in[bdep_j];
					bdep_j = bdep_j + 1;
				end
			end
	end
	wire [62:0] clmul_raw_d;
	assign clmul_raw_d[62:0] = ((((((((((((((((((((((((((((((({63 {rs2_in[0]}} & {31'b0000000000000000000000000000000, rs1_in[31:0]}) ^ ({63 {rs2_in[1]}} & {30'b000000000000000000000000000000, rs1_in[31:0], 1'b0})) ^ ({63 {rs2_in[2]}} & {29'b00000000000000000000000000000, rs1_in[31:0], 2'b00})) ^ ({63 {rs2_in[3]}} & {28'b0000000000000000000000000000, rs1_in[31:0], 3'b000})) ^ ({63 {rs2_in[4]}} & {27'b000000000000000000000000000, rs1_in[31:0], 4'b0000})) ^ ({63 {rs2_in[5]}} & {26'b00000000000000000000000000, rs1_in[31:0], 5'b00000})) ^ ({63 {rs2_in[6]}} & {25'b0000000000000000000000000, rs1_in[31:0], 6'b000000})) ^ ({63 {rs2_in[7]}} & {24'b000000000000000000000000, rs1_in[31:0], 7'b0000000})) ^ ({63 {rs2_in[8]}} & {23'b00000000000000000000000, rs1_in[31:0], 8'b00000000})) ^ ({63 {rs2_in[9]}} & {22'b0000000000000000000000, rs1_in[31:0], 9'b000000000})) ^ ({63 {rs2_in[10]}} & {21'b000000000000000000000, rs1_in[31:0], 10'b0000000000})) ^ ({63 {rs2_in[11]}} & {20'b00000000000000000000, rs1_in[31:0], 11'b00000000000})) ^ ({63 {rs2_in[12]}} & {19'b0000000000000000000, rs1_in[31:0], 12'b000000000000})) ^ ({63 {rs2_in[13]}} & {18'b000000000000000000, rs1_in[31:0], 13'b0000000000000})) ^ ({63 {rs2_in[14]}} & {17'b00000000000000000, rs1_in[31:0], 14'b00000000000000})) ^ ({63 {rs2_in[15]}} & {16'b0000000000000000, rs1_in[31:0], 15'b000000000000000})) ^ ({63 {rs2_in[16]}} & {15'b000000000000000, rs1_in[31:0], 16'b0000000000000000})) ^ ({63 {rs2_in[17]}} & {14'b00000000000000, rs1_in[31:0], 17'b00000000000000000})) ^ ({63 {rs2_in[18]}} & {13'b0000000000000, rs1_in[31:0], 18'b000000000000000000})) ^ ({63 {rs2_in[19]}} & {12'b000000000000, rs1_in[31:0], 19'b0000000000000000000})) ^ ({63 {rs2_in[20]}} & {11'b00000000000, rs1_in[31:0], 20'b00000000000000000000})) ^ ({63 {rs2_in[21]}} & {10'b0000000000, rs1_in[31:0], 21'b000000000000000000000})) ^ ({63 {rs2_in[22]}} & {9'b000000000, rs1_in[31:0], 22'b0000000000000000000000})) ^ ({63 {rs2_in[23]}} & {8'b00000000, rs1_in[31:0], 23'b00000000000000000000000})) ^ ({63 {rs2_in[24]}} & {7'b0000000, rs1_in[31:0], 24'b000000000000000000000000})) ^ ({63 {rs2_in[25]}} & {6'b000000, rs1_in[31:0], 25'b0000000000000000000000000})) ^ ({63 {rs2_in[26]}} & {5'b00000, rs1_in[31:0], 26'b00000000000000000000000000})) ^ ({63 {rs2_in[27]}} & {4'b0000, rs1_in[31:0], 27'b000000000000000000000000000})) ^ ({63 {rs2_in[28]}} & {3'b000, rs1_in[31:0], 28'b0000000000000000000000000000})) ^ ({63 {rs2_in[29]}} & {2'b00, rs1_in[31:0], 29'b00000000000000000000000000000})) ^ ({63 {rs2_in[30]}} & {1'b0, rs1_in[31:0], 30'b000000000000000000000000000000})) ^ ({63 {rs2_in[31]}} & {rs1_in[31:0], 31'b0000000000000000000000000000000});
	wire [31:0] grev1_d;
	wire [31:0] grev2_d;
	wire [31:0] grev4_d;
	wire [31:0] grev8_d;
	wire [31:0] grev_d;
	assign grev1_d[31:0] = (rs2_in[0] ? {rs1_in[30], rs1_in[31], rs1_in[28], rs1_in[29], rs1_in[26], rs1_in[27], rs1_in[24], rs1_in[25], rs1_in[22], rs1_in[23], rs1_in[20], rs1_in[21], rs1_in[18], rs1_in[19], rs1_in[16], rs1_in[17], rs1_in[14], rs1_in[15], rs1_in[12], rs1_in[13], rs1_in[10], rs1_in[11], rs1_in[8], rs1_in[9], rs1_in[6], rs1_in[7], rs1_in[4], rs1_in[5], rs1_in[2], rs1_in[3], rs1_in[0], rs1_in[1]} : rs1_in[31:0]);
	assign grev2_d[31:0] = (rs2_in[1] ? {grev1_d[29:28], grev1_d[31:30], grev1_d[25:24], grev1_d[27:26], grev1_d[21:20], grev1_d[23:22], grev1_d[17:16], grev1_d[19:18], grev1_d[13:12], grev1_d[15:14], grev1_d[9:8], grev1_d[11:10], grev1_d[5:4], grev1_d[7:6], grev1_d[1:0], grev1_d[3:2]} : grev1_d[31:0]);
	assign grev4_d[31:0] = (rs2_in[2] ? {grev2_d[27:24], grev2_d[31:28], grev2_d[19:16], grev2_d[23:20], grev2_d[11:8], grev2_d[15:12], grev2_d[3:0], grev2_d[7:4]} : grev2_d[31:0]);
	assign grev8_d[31:0] = (rs2_in[3] ? {grev4_d[23:16], grev4_d[31:24], grev4_d[7:0], grev4_d[15:8]} : grev4_d[31:0]);
	assign grev_d[31:0] = (rs2_in[4] ? {grev8_d[15:0], grev8_d[31:16]} : grev8_d[31:0]);
	wire [31:0] gorc1_d;
	wire [31:0] gorc2_d;
	wire [31:0] gorc4_d;
	wire [31:0] gorc8_d;
	wire [31:0] gorc_d;
	assign gorc1_d[31:0] = ({32 {rs2_in[0]}} & {rs1_in[30], rs1_in[31], rs1_in[28], rs1_in[29], rs1_in[26], rs1_in[27], rs1_in[24], rs1_in[25], rs1_in[22], rs1_in[23], rs1_in[20], rs1_in[21], rs1_in[18], rs1_in[19], rs1_in[16], rs1_in[17], rs1_in[14], rs1_in[15], rs1_in[12], rs1_in[13], rs1_in[10], rs1_in[11], rs1_in[8], rs1_in[9], rs1_in[6], rs1_in[7], rs1_in[4], rs1_in[5], rs1_in[2], rs1_in[3], rs1_in[0], rs1_in[1]}) | rs1_in[31:0];
	assign gorc2_d[31:0] = ({32 {rs2_in[1]}} & {gorc1_d[29:28], gorc1_d[31:30], gorc1_d[25:24], gorc1_d[27:26], gorc1_d[21:20], gorc1_d[23:22], gorc1_d[17:16], gorc1_d[19:18], gorc1_d[13:12], gorc1_d[15:14], gorc1_d[9:8], gorc1_d[11:10], gorc1_d[5:4], gorc1_d[7:6], gorc1_d[1:0], gorc1_d[3:2]}) | gorc1_d[31:0];
	assign gorc4_d[31:0] = ({32 {rs2_in[2]}} & {gorc2_d[27:24], gorc2_d[31:28], gorc2_d[19:16], gorc2_d[23:20], gorc2_d[11:8], gorc2_d[15:12], gorc2_d[3:0], gorc2_d[7:4]}) | gorc2_d[31:0];
	assign gorc8_d[31:0] = ({32 {rs2_in[3]}} & {gorc4_d[23:16], gorc4_d[31:24], gorc4_d[7:0], gorc4_d[15:8]}) | gorc4_d[31:0];
	assign gorc_d[31:0] = ({32 {rs2_in[4]}} & {gorc8_d[15:0], gorc8_d[31:16]}) | gorc8_d[31:0];
	wire [31:0] shfl8_d;
	wire [31:0] shfl4_d;
	wire [31:0] shfl2_d;
	wire [31:0] shfl_d;
	assign shfl8_d[31:0] = (rs2_in[3] ? {rs1_in[31:24], rs1_in[15:8], rs1_in[23:16], rs1_in[7:0]} : rs1_in[31:0]);
	assign shfl4_d[31:0] = (rs2_in[2] ? {shfl8_d[31:28], shfl8_d[23:20], shfl8_d[27:24], shfl8_d[19:16], shfl8_d[15:12], shfl8_d[7:4], shfl8_d[11:8], shfl8_d[3:0]} : shfl8_d[31:0]);
	assign shfl2_d[31:0] = (rs2_in[1] ? {shfl4_d[31:30], shfl4_d[27:26], shfl4_d[29:28], shfl4_d[25:24], shfl4_d[23:22], shfl4_d[19:18], shfl4_d[21:20], shfl4_d[17:16], shfl4_d[15:14], shfl4_d[11:10], shfl4_d[13:12], shfl4_d[9:8], shfl4_d[7:6], shfl4_d[3:2], shfl4_d[5:4], shfl4_d[1:0]} : shfl4_d[31:0]);
	assign shfl_d[31:0] = (rs2_in[0] ? {shfl2_d[31], shfl2_d[29], shfl2_d[30], shfl2_d[28], shfl2_d[27], shfl2_d[25], shfl2_d[26], shfl2_d[24], shfl2_d[23], shfl2_d[21], shfl2_d[22], shfl2_d[20], shfl2_d[19], shfl2_d[17], shfl2_d[18], shfl2_d[16], shfl2_d[15], shfl2_d[13], shfl2_d[14], shfl2_d[12], shfl2_d[11], shfl2_d[9], shfl2_d[10], shfl2_d[8], shfl2_d[7], shfl2_d[5], shfl2_d[6], shfl2_d[4], shfl2_d[3], shfl2_d[1], shfl2_d[2], shfl2_d[0]} : shfl2_d[31:0]);
	wire [31:0] unshfl1_d;
	wire [31:0] unshfl2_d;
	wire [31:0] unshfl4_d;
	wire [31:0] unshfl_d;
	assign unshfl1_d[31:0] = (rs2_in[0] ? {rs1_in[31], rs1_in[29], rs1_in[30], rs1_in[28], rs1_in[27], rs1_in[25], rs1_in[26], rs1_in[24], rs1_in[23], rs1_in[21], rs1_in[22], rs1_in[20], rs1_in[19], rs1_in[17], rs1_in[18], rs1_in[16], rs1_in[15], rs1_in[13], rs1_in[14], rs1_in[12], rs1_in[11], rs1_in[9], rs1_in[10], rs1_in[8], rs1_in[7], rs1_in[5], rs1_in[6], rs1_in[4], rs1_in[3], rs1_in[1], rs1_in[2], rs1_in[0]} : rs1_in[31:0]);
	assign unshfl2_d[31:0] = (rs2_in[1] ? {unshfl1_d[31:30], unshfl1_d[27:26], unshfl1_d[29:28], unshfl1_d[25:24], unshfl1_d[23:22], unshfl1_d[19:18], unshfl1_d[21:20], unshfl1_d[17:16], unshfl1_d[15:14], unshfl1_d[11:10], unshfl1_d[13:12], unshfl1_d[9:8], unshfl1_d[7:6], unshfl1_d[3:2], unshfl1_d[5:4], unshfl1_d[1:0]} : unshfl1_d[31:0]);
	assign unshfl4_d[31:0] = (rs2_in[2] ? {unshfl2_d[31:28], unshfl2_d[23:20], unshfl2_d[27:24], unshfl2_d[19:16], unshfl2_d[15:12], unshfl2_d[7:4], unshfl2_d[11:8], unshfl2_d[3:0]} : unshfl2_d[31:0]);
	assign unshfl_d[31:0] = (rs2_in[3] ? {unshfl4_d[31:24], unshfl4_d[15:8], unshfl4_d[23:16], unshfl4_d[7:0]} : unshfl4_d[31:0]);
	wire crc32_all;
	wire [31:0] crc32_poly_rev;
	wire [31:0] crc32c_poly_rev;
	integer crc32_bi;
	integer crc32_hi;
	integer crc32_wi;
	integer crc32c_bi;
	integer crc32c_hi;
	integer crc32c_wi;
	reg [31:0] crc32_bd;
	reg [31:0] crc32_hd;
	reg [31:0] crc32_wd;
	reg [31:0] crc32c_bd;
	reg [31:0] crc32c_hd;
	reg [31:0] crc32c_wd;
	assign crc32_all = ((((ap_crc32_b | ap_crc32_h) | ap_crc32_w) | ap_crc32c_b) | ap_crc32c_h) | ap_crc32c_w;
	assign crc32_poly_rev[31:0] = 32'hedb88320;
	assign crc32c_poly_rev[31:0] = 32'h82f63b78;
	always @(*) begin
		crc32_bd[31:0] = rs1_in[31:0];
		for (crc32_bi = 0; crc32_bi < 8; crc32_bi = crc32_bi + 1)
			crc32_bd[31:0] = (crc32_bd[31:0] >> 1) ^ (crc32_poly_rev[31:0] & {32 {crc32_bd[0]}});
	end
	always @(*) begin
		crc32_hd[31:0] = rs1_in[31:0];
		for (crc32_hi = 0; crc32_hi < 16; crc32_hi = crc32_hi + 1)
			crc32_hd[31:0] = (crc32_hd[31:0] >> 1) ^ (crc32_poly_rev[31:0] & {32 {crc32_hd[0]}});
	end
	always @(*) begin
		crc32_wd[31:0] = rs1_in[31:0];
		for (crc32_wi = 0; crc32_wi < 32; crc32_wi = crc32_wi + 1)
			crc32_wd[31:0] = (crc32_wd[31:0] >> 1) ^ (crc32_poly_rev[31:0] & {32 {crc32_wd[0]}});
	end
	always @(*) begin
		crc32c_bd[31:0] = rs1_in[31:0];
		for (crc32c_bi = 0; crc32c_bi < 8; crc32c_bi = crc32c_bi + 1)
			crc32c_bd[31:0] = (crc32c_bd[31:0] >> 1) ^ (crc32c_poly_rev[31:0] & {32 {crc32c_bd[0]}});
	end
	always @(*) begin
		crc32c_hd[31:0] = rs1_in[31:0];
		for (crc32c_hi = 0; crc32c_hi < 16; crc32c_hi = crc32c_hi + 1)
			crc32c_hd[31:0] = (crc32c_hd[31:0] >> 1) ^ (crc32c_poly_rev[31:0] & {32 {crc32c_hd[0]}});
	end
	always @(*) begin
		crc32c_wd[31:0] = rs1_in[31:0];
		for (crc32c_wi = 0; crc32c_wi < 32; crc32c_wi = crc32c_wi + 1)
			crc32c_wd[31:0] = (crc32c_wd[31:0] >> 1) ^ (crc32c_poly_rev[31:0] & {32 {crc32c_wd[0]}});
	end
	wire [4:0] bfp_len;
	wire [4:0] bfp_off;
	wire [31:0] bfp_len_mask_;
	wire [15:0] bfp_preshift_data;
	wire [63:0] bfp_shift_data;
	wire [63:0] bfp_shift_mask;
	wire [31:0] bfp_result_d;
	assign bfp_len[3:0] = rs2_in[27:24];
	assign bfp_len[4] = bfp_len[3:0] == 4'b0000;
	assign bfp_off[4:0] = rs2_in[20:16];
	assign bfp_len_mask_[31:0] = 32'hffffffff << bfp_len[4:0];
	assign bfp_preshift_data[15:0] = rs2_in[15:0] & ~bfp_len_mask_[15:0];
	assign bfp_shift_data[63:0] = {16'b0000000000000000, bfp_preshift_data[15:0], 16'b0000000000000000, bfp_preshift_data[15:0]} << bfp_off[4:0];
	assign bfp_shift_mask[63:0] = {bfp_len_mask_[31:0], bfp_len_mask_[31:0]} << bfp_off[4:0];
	assign bfp_result_d[31:0] = bfp_shift_data[63:32] | (rs1_in[31:0] & bfp_shift_mask[63:32]);
	assign bitmanip_sel_d = (((((((((ap_bext | ap_bdep) | ap_clmul) | ap_clmulh) | ap_clmulr) | ap_grev) | ap_gorc) | ap_shfl) | ap_unshfl) | crc32_all) | ap_bfp;
	assign bitmanip_d[31:0] = ((((((((((((((({32 {ap_bext}} & bext_d[31:0]) | ({32 {ap_bdep}} & bdep_d[31:0])) | ({32 {ap_clmul}} & clmul_raw_d[31:0])) | ({32 {ap_clmulh}} & {1'b0, clmul_raw_d[62:32]})) | ({32 {ap_clmulr}} & clmul_raw_d[62:31])) | ({32 {ap_grev}} & grev_d[31:0])) | ({32 {ap_gorc}} & gorc_d[31:0])) | ({32 {ap_shfl}} & shfl_d[31:0])) | ({32 {ap_unshfl}} & unshfl_d[31:0])) | ({32 {ap_crc32_b}} & crc32_bd[31:0])) | ({32 {ap_crc32_h}} & crc32_hd[31:0])) | ({32 {ap_crc32_w}} & crc32_wd[31:0])) | ({32 {ap_crc32c_b}} & crc32c_bd[31:0])) | ({32 {ap_crc32c_h}} & crc32c_hd[31:0])) | ({32 {ap_crc32c_w}} & crc32c_wd[31:0])) | ({32 {ap_bfp}} & bfp_result_d[31:0]);
	rvdffe #(.WIDTH(33)) i_bitmanip_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din({bitmanip_sel_d, bitmanip_d[31:0]}),
		.dout({bitmanip_sel_x, bitmanip_x[31:0]}),
		.en(bit_x_enable)
	);
	assign result_x[31:0] = (({32 {~bitmanip_sel_x & ~low_x}} & prod_x[63:32]) | ({32 {~bitmanip_sel_x & low_x}} & prod_x[31:0])) | bitmanip_x[31:0];
endmodule
module eb1_ifu (
	free_l2clk,
	active_clk,
	clk,
	rst_l,
	dec_i0_decode_d,
	exu_flush_final,
	dec_tlu_i0_commit_cmt,
	dec_tlu_flush_err_wb,
	dec_tlu_flush_noredir_wb,
	exu_flush_path_final,
	dec_tlu_mrac_ff,
	dec_tlu_fence_i_wb,
	dec_tlu_flush_leak_one_wb,
	dec_tlu_bpred_disable,
	dec_tlu_core_ecc_disable,
	dec_tlu_force_halt,
	ifu_axi_awvalid,
	ifu_axi_awid,
	ifu_axi_awaddr,
	ifu_axi_awregion,
	ifu_axi_awlen,
	ifu_axi_awsize,
	ifu_axi_awburst,
	ifu_axi_awlock,
	ifu_axi_awcache,
	ifu_axi_awprot,
	ifu_axi_awqos,
	ifu_axi_wvalid,
	ifu_axi_wdata,
	ifu_axi_wstrb,
	ifu_axi_wlast,
	ifu_axi_bready,
	ifu_axi_arvalid,
	ifu_axi_arready,
	ifu_axi_arid,
	ifu_axi_araddr,
	ifu_axi_arregion,
	ifu_axi_arlen,
	ifu_axi_arsize,
	ifu_axi_arburst,
	ifu_axi_arlock,
	ifu_axi_arcache,
	ifu_axi_arprot,
	ifu_axi_arqos,
	ifu_axi_rvalid,
	ifu_axi_rready,
	ifu_axi_rid,
	ifu_axi_rdata,
	ifu_axi_rresp,
	ifu_bus_clk_en,
	dma_iccm_req,
	dma_mem_addr,
	dma_mem_sz,
	dma_mem_write,
	dma_mem_wdata,
	dma_mem_tag,
	dma_iccm_stall_any,
	iccm_dma_ecc_error,
	iccm_dma_rvalid,
	iccm_dma_rdata,
	iccm_dma_rtag,
	iccm_ready,
	ifu_pmu_instr_aligned,
	ifu_pmu_fetch_stall,
	ifu_ic_error_start,
	ic_rw_addr,
	ic_wr_en,
	ic_rd_en,
	ic_wr_data,
	ic_rd_data,
	ic_debug_rd_data,
	ictag_debug_rd_data,
	ic_debug_wr_data,
	ifu_ic_debug_rd_data,
	ic_eccerr,
	ic_parerr,
	ic_premux_data,
	ic_sel_premux_data,
	ic_debug_addr,
	ic_debug_rd_en,
	ic_debug_wr_en,
	ic_debug_tag_array,
	ic_debug_way,
	ic_tag_valid,
	ic_rd_hit,
	ic_tag_perr,
	iccm_rw_addr,
	iccm_wren,
	iccm_rden,
	iccm_wr_data,
	iccm_wr_size,
	iccm_rd_data,
	iccm_rd_data_ecc,
	ifu_iccm_rd_ecc_single_err,
	ifu_pmu_ic_miss,
	ifu_pmu_ic_hit,
	ifu_pmu_bus_error,
	ifu_pmu_bus_busy,
	ifu_pmu_bus_trxn,
	ifu_i0_icaf,
	ifu_i0_icaf_type,
	ifu_i0_valid,
	ifu_i0_icaf_second,
	ifu_i0_dbecc,
	iccm_dma_sb_error,
	ifu_i0_instr,
	ifu_i0_pc,
	ifu_i0_pc4,
	ifu_miss_state_idle,
	i0_brp,
	ifu_i0_bp_index,
	ifu_i0_bp_fghr,
	ifu_i0_bp_btag,
	ifu_i0_fa_index,
	exu_mp_pkt,
	exu_mp_eghr,
	exu_mp_fghr,
	exu_mp_index,
	exu_mp_btag,
	dec_tlu_br0_r_pkt,
	exu_i0_br_fghr_r,
	exu_i0_br_index_r,
	dec_fa_error_index,
	dec_tlu_flush_lower_wb,
	ifu_i0_cinst,
	dec_tlu_ic_diag_pkt,
	ifu_ic_debug_rd_data_valid,
	iccm_buf_correct_ecc,
	iccm_correction_state,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire free_l2clk;
	input wire active_clk;
	input wire clk;
	input wire rst_l;
	input wire dec_i0_decode_d;
	input wire exu_flush_final;
	input wire dec_tlu_i0_commit_cmt;
	input wire dec_tlu_flush_err_wb;
	input wire dec_tlu_flush_noredir_wb;
	input wire [31:1] exu_flush_path_final;
	input wire [31:0] dec_tlu_mrac_ff;
	input wire dec_tlu_fence_i_wb;
	input wire dec_tlu_flush_leak_one_wb;
	input wire dec_tlu_bpred_disable;
	input wire dec_tlu_core_ecc_disable;
	input wire dec_tlu_force_halt;
	output wire ifu_axi_awvalid;
	output wire [pt[826-:8] - 1:0] ifu_axi_awid;
	output wire [31:0] ifu_axi_awaddr;
	output wire [3:0] ifu_axi_awregion;
	output wire [7:0] ifu_axi_awlen;
	output wire [2:0] ifu_axi_awsize;
	output wire [1:0] ifu_axi_awburst;
	output wire ifu_axi_awlock;
	output wire [3:0] ifu_axi_awcache;
	output wire [2:0] ifu_axi_awprot;
	output wire [3:0] ifu_axi_awqos;
	output wire ifu_axi_wvalid;
	output wire [63:0] ifu_axi_wdata;
	output wire [7:0] ifu_axi_wstrb;
	output wire ifu_axi_wlast;
	output wire ifu_axi_bready;
	output wire ifu_axi_arvalid;
	input wire ifu_axi_arready;
	output wire [pt[826-:8] - 1:0] ifu_axi_arid;
	output wire [31:0] ifu_axi_araddr;
	output wire [3:0] ifu_axi_arregion;
	output wire [7:0] ifu_axi_arlen;
	output wire [2:0] ifu_axi_arsize;
	output wire [1:0] ifu_axi_arburst;
	output wire ifu_axi_arlock;
	output wire [3:0] ifu_axi_arcache;
	output wire [2:0] ifu_axi_arprot;
	output wire [3:0] ifu_axi_arqos;
	input wire ifu_axi_rvalid;
	output wire ifu_axi_rready;
	input wire [pt[826-:8] - 1:0] ifu_axi_rid;
	input wire [63:0] ifu_axi_rdata;
	input wire [1:0] ifu_axi_rresp;
	input wire ifu_bus_clk_en;
	input wire dma_iccm_req;
	input wire [31:0] dma_mem_addr;
	input wire [2:0] dma_mem_sz;
	input wire dma_mem_write;
	input wire [63:0] dma_mem_wdata;
	input wire [2:0] dma_mem_tag;
	input wire dma_iccm_stall_any;
	output wire iccm_dma_ecc_error;
	output wire iccm_dma_rvalid;
	output wire [63:0] iccm_dma_rdata;
	output wire [2:0] iccm_dma_rtag;
	output wire iccm_ready;
	output wire ifu_pmu_instr_aligned;
	output wire ifu_pmu_fetch_stall;
	output wire ifu_ic_error_start;
	output wire [31:1] ic_rw_addr;
	output wire [pt[1060-:7] - 1:0] ic_wr_en;
	output wire ic_rd_en;
	output wire [(pt[1189-:7] * 71) - 1:0] ic_wr_data;
	input wire [63:0] ic_rd_data;
	input wire [70:0] ic_debug_rd_data;
	input wire [25:0] ictag_debug_rd_data;
	output wire [70:0] ic_debug_wr_data;
	output wire [70:0] ifu_ic_debug_rd_data;
	input wire [pt[1189-:7] - 1:0] ic_eccerr;
	input wire [pt[1189-:7] - 1:0] ic_parerr;
	output wire [63:0] ic_premux_data;
	output wire ic_sel_premux_data;
	output wire [pt[1104-:9]:3] ic_debug_addr;
	output wire ic_debug_rd_en;
	output wire ic_debug_wr_en;
	output wire ic_debug_tag_array;
	output wire [pt[1060-:7] - 1:0] ic_debug_way;
	output wire [pt[1060-:7] - 1:0] ic_tag_valid;
	input wire [pt[1060-:7] - 1:0] ic_rd_hit;
	input wire ic_tag_perr;
	output wire [pt[936-:9] - 1:1] iccm_rw_addr;
	output wire iccm_wren;
	output wire iccm_rden;
	output wire [77:0] iccm_wr_data;
	output wire [2:0] iccm_wr_size;
	input wire [63:0] iccm_rd_data;
	input wire [77:0] iccm_rd_data_ecc;
	output wire ifu_iccm_rd_ecc_single_err;
	output wire ifu_pmu_ic_miss;
	output wire ifu_pmu_ic_hit;
	output wire ifu_pmu_bus_error;
	output wire ifu_pmu_bus_busy;
	output wire ifu_pmu_bus_trxn;
	output wire ifu_i0_icaf;
	output wire [1:0] ifu_i0_icaf_type;
	output wire ifu_i0_valid;
	output wire ifu_i0_icaf_second;
	output wire ifu_i0_dbecc;
	output wire iccm_dma_sb_error;
	output wire [31:0] ifu_i0_instr;
	output wire [31:1] ifu_i0_pc;
	output wire ifu_i0_pc4;
	output wire ifu_miss_state_idle;
	output wire [50:0] i0_brp;
	output wire [pt[2172-:9]:pt[2163-:6]] ifu_i0_bp_index;
	output wire [pt[2236-:8] - 1:0] ifu_i0_bp_fghr;
	output wire [pt[2139-:9] - 1:0] ifu_i0_bp_btag;
	output wire [$clog2(pt[2061-:14]) - 1:0] ifu_i0_fa_index;
	input wire [55:0] exu_mp_pkt;
	input wire [pt[2236-:8] - 1:0] exu_mp_eghr;
	input wire [pt[2236-:8] - 1:0] exu_mp_fghr;
	input wire [pt[2172-:9]:pt[2163-:6]] exu_mp_index;
	input wire [pt[2139-:9] - 1:0] exu_mp_btag;
	input wire [6:0] dec_tlu_br0_r_pkt;
	input wire [pt[2236-:8] - 1:0] exu_i0_br_fghr_r;
	input wire [pt[2172-:9]:pt[2163-:6]] exu_i0_br_index_r;
	input wire [$clog2(pt[2061-:14]) - 1:0] dec_fa_error_index;
	input dec_tlu_flush_lower_wb;
	output wire [15:0] ifu_i0_cinst;
	input wire [89:0] dec_tlu_ic_diag_pkt;
	output wire ifu_ic_debug_rd_data_valid;
	output wire iccm_buf_correct_ecc;
	output wire iccm_correction_state;
	input wire scan_mode;
	localparam TAGWIDTH = 2;
	localparam IDWIDTH = 2;
	wire ifu_fb_consume1;
	wire ifu_fb_consume2;
	wire [31:1] ifc_fetch_addr_f;
	wire [31:1] ifc_fetch_addr_bf;
	wire [1:0] ifu_fetch_val;
	wire [31:1] ifu_fetch_pc;
	wire iccm_rd_ecc_single_err;
	wire ic_error_start;
	assign ifu_iccm_rd_ecc_single_err = iccm_rd_ecc_single_err;
	assign ifu_ic_error_start = ic_error_start;
	wire ic_write_stall;
	wire ic_dma_active;
	wire ifc_dma_access_ok;
	wire [1:0] ic_access_fault_f;
	wire [1:0] ic_access_fault_type_f;
	wire ifu_ic_mb_empty;
	wire ic_hit_f;
	wire [1:0] ifu_bp_way_f;
	wire ifu_bp_hit_taken_f;
	wire [31:1] ifu_bp_btb_target_f;
	wire ifu_bp_inst_mask_f;
	wire [1:0] ifu_bp_hist1_f;
	wire [1:0] ifu_bp_hist0_f;
	wire [11:0] ifu_bp_poffset_f;
	wire [1:0] ifu_bp_ret_f;
	wire [1:0] ifu_bp_pc4_f;
	wire [1:0] ifu_bp_valid_f;
	wire [pt[2236-:8] - 1:0] ifu_bp_fghr_f;
	wire [(2 * $clog2(pt[2061-:14])) - 1:0] ifu_bp_fa_index_f;
	wire ifc_fetch_req_bf;
	wire ifc_fetch_req_bf_raw;
	wire ifc_fetch_req_f;
	wire ifc_fetch_uncacheable_bf;
	wire ifc_iccm_access_bf;
	wire ifc_region_acc_fault_bf;
	eb1_ifu_ifc_ctl #(.pt(pt)) ifc(
		.clk(clk),
		.free_l2clk(free_l2clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.ic_hit_f(ic_hit_f),
		.ifu_ic_mb_empty(ifu_ic_mb_empty),
		.ifu_fb_consume1(ifu_fb_consume1),
		.ifu_fb_consume2(ifu_fb_consume2),
		.dec_tlu_flush_noredir_wb(dec_tlu_flush_noredir_wb),
		.exu_flush_final(exu_flush_final),
		.exu_flush_path_final(exu_flush_path_final),
		.ifu_bp_hit_taken_f(ifu_bp_hit_taken_f),
		.ifu_bp_btb_target_f(ifu_bp_btb_target_f),
		.ic_dma_active(ic_dma_active),
		.ic_write_stall(ic_write_stall),
		.dma_iccm_stall_any(dma_iccm_stall_any),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.ifc_fetch_addr_f(ifc_fetch_addr_f),
		.ifc_fetch_addr_bf(ifc_fetch_addr_bf),
		.ifc_fetch_req_f(ifc_fetch_req_f),
		.ifu_pmu_fetch_stall(ifu_pmu_fetch_stall),
		.ifc_fetch_uncacheable_bf(ifc_fetch_uncacheable_bf),
		.ifc_fetch_req_bf(ifc_fetch_req_bf),
		.ifc_fetch_req_bf_raw(ifc_fetch_req_bf_raw),
		.ifc_iccm_access_bf(ifc_iccm_access_bf),
		.ifc_region_acc_fault_bf(ifc_region_acc_fault_bf),
		.ifc_dma_access_ok(ifc_dma_access_ok)
	);
	generate
		if (pt[2130-:5] == 1) begin : bpred
			eb1_ifu_bp_ctl #(.pt(pt)) bp(
				.clk(clk),
				.rst_l(rst_l),
				.ic_hit_f(ic_hit_f),
				.ifc_fetch_addr_f(ifc_fetch_addr_f),
				.ifc_fetch_req_f(ifc_fetch_req_f),
				.dec_tlu_br0_r_pkt(dec_tlu_br0_r_pkt),
				.exu_i0_br_fghr_r(exu_i0_br_fghr_r),
				.exu_i0_br_index_r(exu_i0_br_index_r),
				.dec_fa_error_index(dec_fa_error_index),
				.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_wb),
				.dec_tlu_flush_leak_one_wb(dec_tlu_flush_leak_one_wb),
				.dec_tlu_bpred_disable(dec_tlu_bpred_disable),
				.exu_mp_pkt(exu_mp_pkt),
				.exu_mp_eghr(exu_mp_eghr),
				.exu_mp_fghr(exu_mp_fghr),
				.exu_mp_index(exu_mp_index),
				.exu_mp_btag(exu_mp_btag),
				.exu_flush_final(exu_flush_final),
				.ifu_bp_hit_taken_f(ifu_bp_hit_taken_f),
				.ifu_bp_btb_target_f(ifu_bp_btb_target_f),
				.ifu_bp_inst_mask_f(ifu_bp_inst_mask_f),
				.ifu_bp_fghr_f(ifu_bp_fghr_f),
				.ifu_bp_way_f(ifu_bp_way_f),
				.ifu_bp_ret_f(ifu_bp_ret_f),
				.ifu_bp_hist1_f(ifu_bp_hist1_f),
				.ifu_bp_hist0_f(ifu_bp_hist0_f),
				.ifu_bp_pc4_f(ifu_bp_pc4_f),
				.ifu_bp_valid_f(ifu_bp_valid_f),
				.ifu_bp_poffset_f(ifu_bp_poffset_f),
				.ifu_bp_fa_index_f(ifu_bp_fa_index_f),
				.scan_mode(scan_mode)
			);
		end
		else begin : bpred
			assign ifu_bp_hit_taken_f = 1'b0;
			wire btb_wr_en_way0;
			wire btb_wr_en_way1;
			wire dec_tlu_error_wb;
			wire [16 + pt[2139-:9]:0] btb_wr_data;
			assign btb_wr_en_way0 = 1'b0;
			assign btb_wr_en_way1 = 1'b0;
			assign btb_wr_data = {((16 + pt[2139-:9]) >= 0 ? (16 + pt[2139-:9]) + 1 : 1 - (16 + pt[2139-:9])) {1'sb0}};
			assign dec_tlu_error_wb = 1'b0;
			assign ifu_bp_inst_mask_f = 1'b1;
		end
	endgenerate
	wire [1:0] ic_fetch_val_f;
	wire [31:0] ic_data_f;
	wire [31:0] ifu_fetch_data_f;
	wire ifc_fetch_req_f_raw;
	wire [1:0] iccm_rd_ecc_double_err;
	wire ifu_async_error_start;
	assign ifu_fetch_data_f[31:0] = ic_data_f[31:0];
	assign ifu_fetch_val[1:0] = ic_fetch_val_f[1:0];
	assign ifu_fetch_pc[31:1] = ifc_fetch_addr_f[31:1];
	eb1_ifu_aln_ctl #(.pt(pt)) aln(
		.scan_mode(scan_mode),
		.rst_l(rst_l),
		.clk(clk),
		.active_clk(active_clk),
		.ifu_async_error_start(ifu_async_error_start),
		.iccm_rd_ecc_double_err(iccm_rd_ecc_double_err),
		.ic_access_fault_f(ic_access_fault_f),
		.ic_access_fault_type_f(ic_access_fault_type_f),
		.exu_flush_final(exu_flush_final),
		.dec_i0_decode_d(dec_i0_decode_d),
		.ifu_fetch_data_f(ifu_fetch_data_f),
		.ifu_fetch_val(ifu_fetch_val),
		.ifu_fetch_pc(ifu_fetch_pc),
		.ifu_i0_valid(ifu_i0_valid),
		.ifu_i0_icaf(ifu_i0_icaf),
		.ifu_i0_icaf_type(ifu_i0_icaf_type),
		.ifu_i0_icaf_second(ifu_i0_icaf_second),
		.ifu_i0_dbecc(ifu_i0_dbecc),
		.ifu_i0_instr(ifu_i0_instr),
		.ifu_i0_pc(ifu_i0_pc),
		.ifu_i0_pc4(ifu_i0_pc4),
		.ifu_fb_consume1(ifu_fb_consume1),
		.ifu_fb_consume2(ifu_fb_consume2),
		.ifu_bp_fghr_f(ifu_bp_fghr_f),
		.ifu_bp_btb_target_f(ifu_bp_btb_target_f),
		.ifu_bp_poffset_f(ifu_bp_poffset_f),
		.ifu_bp_fa_index_f(ifu_bp_fa_index_f),
		.ifu_bp_hist0_f(ifu_bp_hist0_f),
		.ifu_bp_hist1_f(ifu_bp_hist1_f),
		.ifu_bp_pc4_f(ifu_bp_pc4_f),
		.ifu_bp_way_f(ifu_bp_way_f),
		.ifu_bp_valid_f(ifu_bp_valid_f),
		.ifu_bp_ret_f(ifu_bp_ret_f),
		.i0_brp(i0_brp),
		.ifu_i0_bp_index(ifu_i0_bp_index),
		.ifu_i0_bp_fghr(ifu_i0_bp_fghr),
		.ifu_i0_bp_btag(ifu_i0_bp_btag),
		.ifu_i0_fa_index(ifu_i0_fa_index),
		.ifu_pmu_instr_aligned(ifu_pmu_instr_aligned),
		.ifu_i0_cinst(ifu_i0_cinst)
	);
	eb1_ifu_mem_ctl #(.pt(pt)) mem_ctl(
		.clk(clk),
		.active_clk(active_clk),
		.free_l2clk(free_l2clk),
		.rst_l(rst_l),
		.exu_flush_final(exu_flush_final),
		.dec_tlu_flush_lower_wb(dec_tlu_flush_lower_wb),
		.dec_tlu_flush_err_wb(dec_tlu_flush_err_wb),
		.dec_tlu_i0_commit_cmt(dec_tlu_i0_commit_cmt),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.ifc_fetch_addr_bf(ifc_fetch_addr_bf),
		.ifc_fetch_uncacheable_bf(ifc_fetch_uncacheable_bf),
		.ifc_fetch_req_bf(ifc_fetch_req_bf),
		.ifc_fetch_req_bf_raw(ifc_fetch_req_bf_raw),
		.ifc_iccm_access_bf(ifc_iccm_access_bf),
		.ifc_region_acc_fault_bf(ifc_region_acc_fault_bf),
		.ifc_dma_access_ok(ifc_dma_access_ok),
		.dec_tlu_fence_i_wb(dec_tlu_fence_i_wb),
		.ifu_bp_hit_taken_f(ifu_bp_hit_taken_f),
		.ifu_bp_inst_mask_f(ifu_bp_inst_mask_f),
		.ifu_miss_state_idle(ifu_miss_state_idle),
		.ifu_ic_mb_empty(ifu_ic_mb_empty),
		.ic_dma_active(ic_dma_active),
		.ic_write_stall(ic_write_stall),
		.ifu_pmu_ic_miss(ifu_pmu_ic_miss),
		.ifu_pmu_ic_hit(ifu_pmu_ic_hit),
		.ifu_pmu_bus_error(ifu_pmu_bus_error),
		.ifu_pmu_bus_busy(ifu_pmu_bus_busy),
		.ifu_pmu_bus_trxn(ifu_pmu_bus_trxn),
		.ifu_axi_awvalid(ifu_axi_awvalid),
		.ifu_axi_awid(ifu_axi_awid),
		.ifu_axi_awaddr(ifu_axi_awaddr),
		.ifu_axi_awregion(ifu_axi_awregion),
		.ifu_axi_awlen(ifu_axi_awlen),
		.ifu_axi_awsize(ifu_axi_awsize),
		.ifu_axi_awburst(ifu_axi_awburst),
		.ifu_axi_awlock(ifu_axi_awlock),
		.ifu_axi_awcache(ifu_axi_awcache),
		.ifu_axi_awprot(ifu_axi_awprot),
		.ifu_axi_awqos(ifu_axi_awqos),
		.ifu_axi_wvalid(ifu_axi_wvalid),
		.ifu_axi_wdata(ifu_axi_wdata),
		.ifu_axi_wstrb(ifu_axi_wstrb),
		.ifu_axi_wlast(ifu_axi_wlast),
		.ifu_axi_bready(ifu_axi_bready),
		.ifu_axi_arvalid(ifu_axi_arvalid),
		.ifu_axi_arready(ifu_axi_arready),
		.ifu_axi_arid(ifu_axi_arid),
		.ifu_axi_araddr(ifu_axi_araddr),
		.ifu_axi_arregion(ifu_axi_arregion),
		.ifu_axi_arlen(ifu_axi_arlen),
		.ifu_axi_arsize(ifu_axi_arsize),
		.ifu_axi_arburst(ifu_axi_arburst),
		.ifu_axi_arlock(ifu_axi_arlock),
		.ifu_axi_arcache(ifu_axi_arcache),
		.ifu_axi_arprot(ifu_axi_arprot),
		.ifu_axi_arqos(ifu_axi_arqos),
		.ifu_axi_rvalid(ifu_axi_rvalid),
		.ifu_axi_rready(ifu_axi_rready),
		.ifu_axi_rid(ifu_axi_rid),
		.ifu_axi_rdata(ifu_axi_rdata),
		.ifu_axi_rresp(ifu_axi_rresp),
		.ifu_bus_clk_en(ifu_bus_clk_en),
		.dma_iccm_req(dma_iccm_req),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_sz(dma_mem_sz),
		.dma_mem_write(dma_mem_write),
		.dma_mem_wdata(dma_mem_wdata),
		.dma_mem_tag(dma_mem_tag),
		.iccm_dma_ecc_error(iccm_dma_ecc_error),
		.iccm_dma_rvalid(iccm_dma_rvalid),
		.iccm_dma_rdata(iccm_dma_rdata),
		.iccm_dma_rtag(iccm_dma_rtag),
		.iccm_ready(iccm_ready),
		.ic_rw_addr(ic_rw_addr),
		.ic_wr_en(ic_wr_en),
		.ic_rd_en(ic_rd_en),
		.ic_wr_data(ic_wr_data),
		.ic_rd_data(ic_rd_data),
		.ic_debug_rd_data(ic_debug_rd_data),
		.ictag_debug_rd_data(ictag_debug_rd_data),
		.ic_debug_wr_data(ic_debug_wr_data),
		.ifu_ic_debug_rd_data(ifu_ic_debug_rd_data),
		.ic_eccerr(ic_eccerr),
		.ic_parerr(ic_parerr),
		.ic_debug_addr(ic_debug_addr),
		.ic_debug_rd_en(ic_debug_rd_en),
		.ic_debug_wr_en(ic_debug_wr_en),
		.ic_debug_tag_array(ic_debug_tag_array),
		.ic_debug_way(ic_debug_way),
		.ic_tag_valid(ic_tag_valid),
		.ic_rd_hit(ic_rd_hit),
		.ic_tag_perr(ic_tag_perr),
		.iccm_rw_addr(iccm_rw_addr),
		.iccm_wren(iccm_wren),
		.iccm_rden(iccm_rden),
		.iccm_wr_data(iccm_wr_data),
		.iccm_wr_size(iccm_wr_size),
		.iccm_rd_data(iccm_rd_data),
		.iccm_rd_data_ecc(iccm_rd_data_ecc),
		.ifu_fetch_val(ifu_fetch_val),
		.ic_hit_f(ic_hit_f),
		.ic_access_fault_f(ic_access_fault_f),
		.ic_access_fault_type_f(ic_access_fault_type_f),
		.iccm_rd_ecc_single_err(iccm_rd_ecc_single_err),
		.iccm_rd_ecc_double_err(iccm_rd_ecc_double_err),
		.ic_error_start(ic_error_start),
		.ifu_async_error_start(ifu_async_error_start),
		.iccm_dma_sb_error(iccm_dma_sb_error),
		.ic_fetch_val_f(ic_fetch_val_f),
		.ic_premux_data(ic_premux_data),
		.ic_sel_premux_data(ic_sel_premux_data),
		.dec_tlu_ic_diag_pkt(dec_tlu_ic_diag_pkt),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.ifu_ic_debug_rd_data_valid(ifu_ic_debug_rd_data_valid),
		.iccm_buf_correct_ecc(iccm_buf_correct_ecc),
		.iccm_correction_state(iccm_correction_state),
		.scan_mode(scan_mode),
		.ic_data_f(ic_data_f[31:0])
	);
endmodule
module eb1_ifu_aln_ctl (
	scan_mode,
	rst_l,
	clk,
	active_clk,
	ifu_async_error_start,
	iccm_rd_ecc_double_err,
	ic_access_fault_f,
	ic_access_fault_type_f,
	exu_flush_final,
	dec_i0_decode_d,
	ifu_fetch_data_f,
	ifu_fetch_val,
	ifu_fetch_pc,
	ifu_i0_valid,
	ifu_i0_icaf,
	ifu_i0_icaf_type,
	ifu_i0_icaf_second,
	ifu_i0_dbecc,
	ifu_i0_instr,
	ifu_i0_pc,
	ifu_i0_pc4,
	ifu_fb_consume1,
	ifu_fb_consume2,
	ifu_bp_fghr_f,
	ifu_bp_btb_target_f,
	ifu_bp_poffset_f,
	ifu_bp_fa_index_f,
	ifu_bp_hist0_f,
	ifu_bp_hist1_f,
	ifu_bp_pc4_f,
	ifu_bp_way_f,
	ifu_bp_valid_f,
	ifu_bp_ret_f,
	i0_brp,
	ifu_i0_bp_index,
	ifu_i0_bp_fghr,
	ifu_i0_bp_btag,
	ifu_i0_fa_index,
	ifu_pmu_instr_aligned,
	ifu_i0_cinst
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire scan_mode;
	input wire rst_l;
	input wire clk;
	input wire active_clk;
	input wire ifu_async_error_start;
	input wire [1:0] iccm_rd_ecc_double_err;
	input wire [1:0] ic_access_fault_f;
	input wire [1:0] ic_access_fault_type_f;
	input wire exu_flush_final;
	input wire dec_i0_decode_d;
	input wire [31:0] ifu_fetch_data_f;
	input wire [1:0] ifu_fetch_val;
	input wire [31:1] ifu_fetch_pc;
	output wire ifu_i0_valid;
	output wire ifu_i0_icaf;
	output wire [1:0] ifu_i0_icaf_type;
	output wire ifu_i0_icaf_second;
	output wire ifu_i0_dbecc;
	output wire [31:0] ifu_i0_instr;
	output wire [31:1] ifu_i0_pc;
	output wire ifu_i0_pc4;
	output wire ifu_fb_consume1;
	output wire ifu_fb_consume2;
	input wire [pt[2236-:8] - 1:0] ifu_bp_fghr_f;
	input wire [31:1] ifu_bp_btb_target_f;
	input wire [11:0] ifu_bp_poffset_f;
	input wire [(2 * $clog2(pt[2061-:14])) - 1:0] ifu_bp_fa_index_f;
	input wire [1:0] ifu_bp_hist0_f;
	input wire [1:0] ifu_bp_hist1_f;
	input wire [1:0] ifu_bp_pc4_f;
	input wire [1:0] ifu_bp_way_f;
	input wire [1:0] ifu_bp_valid_f;
	input wire [1:0] ifu_bp_ret_f;
	output reg [50:0] i0_brp;
	output wire [pt[2172-:9]:pt[2163-:6]] ifu_i0_bp_index;
	output wire [pt[2236-:8] - 1:0] ifu_i0_bp_fghr;
	output wire [pt[2139-:9] - 1:0] ifu_i0_bp_btag;
	output reg [$clog2(pt[2061-:14]) - 1:0] ifu_i0_fa_index;
	output wire ifu_pmu_instr_aligned;
	output wire [15:0] ifu_i0_cinst;
	wire ifvalid;
	wire shift_f1_f0;
	wire shift_f2_f0;
	wire shift_f2_f1;
	wire fetch_to_f0;
	wire fetch_to_f1;
	wire fetch_to_f2;
	wire [1:0] f2val_in;
	wire [1:0] f2val;
	wire [1:0] f1val_in;
	wire [1:0] f1val;
	wire [1:0] f0val_in;
	wire [1:0] f0val;
	wire [1:0] sf1val;
	wire [1:0] sf0val;
	wire [31:0] aligndata;
	wire first4B;
	wire first2B;
	wire [31:0] uncompress0;
	wire i0_shift;
	wire shift_2B;
	wire shift_4B;
	wire f1_shift_2B;
	wire f2_valid;
	wire sf1_valid;
	wire sf0_valid;
	wire [31:0] ifirst;
	wire [1:0] alignval;
	wire [31:1] firstpc;
	wire [31:1] secondpc;
	wire [11:0] f1poffset;
	wire [11:0] f0poffset;
	wire [pt[2236-:8] - 1:0] f1fghr;
	wire [pt[2236-:8] - 1:0] f0fghr;
	wire [1:0] f1hist1;
	wire [1:0] f0hist1;
	wire [1:0] f1hist0;
	wire [1:0] f0hist0;
	wire [(2 * $clog2(pt[2061-:14])) - 1:0] f0index;
	wire [(2 * $clog2(pt[2061-:14])) - 1:0] f1index;
	wire [(2 * $clog2(pt[2061-:14])) - 1:0] alignindex;
	wire [1:0] f1ictype;
	wire [1:0] f0ictype;
	wire [1:0] f1pc4;
	wire [1:0] f0pc4;
	wire [1:0] f1ret;
	wire [1:0] f0ret;
	wire [1:0] f1way;
	wire [1:0] f0way;
	wire [1:0] f1brend;
	wire [1:0] f0brend;
	wire [1:0] alignbrend;
	wire [1:0] alignpc4;
	wire [1:0] alignret;
	wire [1:0] alignway;
	wire [1:0] alignhist1;
	wire [1:0] alignhist0;
	wire [1:1] alignfromf1;
	reg i0_ends_f1;
	reg i0_br_start_error;
	wire [31:1] f1prett;
	wire [31:1] f0prett;
	wire [1:0] f1dbecc;
	wire [1:0] f0dbecc;
	wire [1:0] f1icaf;
	wire [1:0] f0icaf;
	wire [1:0] aligndbecc;
	wire [1:0] alignicaf;
	reg i0_brp_pc4;
	wire [pt[2172-:9]:pt[2163-:6]] firstpc_hash;
	wire [pt[2172-:9]:pt[2163-:6]] secondpc_hash;
	wire first_legal;
	wire [1:0] wrptr;
	wire [1:0] wrptr_in;
	wire [1:0] rdptr;
	wire [1:0] rdptr_in;
	wire [2:0] qwen;
	wire [31:0] q2;
	wire [31:0] q1;
	wire [31:0] q0;
	wire q2off_in;
	wire q2off;
	wire q1off_in;
	wire q1off;
	wire q0off_in;
	wire q0off;
	wire f0_shift_2B;
	wire [31:0] q0eff;
	wire [31:0] q0final;
	wire q0ptr;
	wire [1:0] q0sel;
	wire [31:0] q1eff;
	wire [15:0] q1final;
	wire q1ptr;
	wire [1:0] q1sel;
	wire [2:0] qren;
	wire consume_fb1;
	wire consume_fb0;
	wire [1:0] icaf_eff;
	localparam BRDATA_SIZE = (pt[2130-:5] ? 16 + (($clog2(pt[2061-:14]) * 2) * pt[2120-:5]) : 2);
	localparam BRDATA_WIDTH = (pt[2130-:5] ? 8 + ($clog2(pt[2061-:14]) * pt[2120-:5]) : 1);
	wire [BRDATA_SIZE - 1:0] brdata_in;
	wire [BRDATA_SIZE - 1:0] brdata2;
	wire [BRDATA_SIZE - 1:0] brdata1;
	wire [BRDATA_SIZE - 1:0] brdata0;
	wire [BRDATA_SIZE - 1:0] brdata1eff;
	wire [BRDATA_SIZE - 1:0] brdata0eff;
	wire [BRDATA_SIZE - 1:0] brdata1final;
	wire [BRDATA_SIZE - 1:0] brdata0final;
	localparam MHI = 1 + (pt[2130-:5] * (43 + pt[2236-:8]));
	localparam MSIZE = 2 + (pt[2130-:5] * (43 + pt[2236-:8]));
	wire [MHI:0] misc_data_in;
	wire [MHI:0] misc2;
	wire [MHI:0] misc1;
	wire [MHI:0] misc0;
	wire [MHI:0] misc1eff;
	wire [MHI:0] misc0eff;
	wire [pt[2139-:9] - 1:0] firstbrtag_hash;
	wire [pt[2139-:9] - 1:0] secondbrtag_hash;
	wire error_stall_in;
	wire error_stall;
	assign error_stall_in = (error_stall | ifu_async_error_start) & ~exu_flush_final;
	rvdff #(.WIDTH(7)) bundle1ff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din({wrptr_in[1:0], rdptr_in[1:0], q2off_in, q1off_in, q0off_in}),
		.dout({wrptr[1:0], rdptr[1:0], q2off, q1off, q0off})
	);
	rvdffie #(
		.WIDTH(7),
		.OVERRIDE(1)
	) bundle2ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din({error_stall_in, f2val_in[1:0], f1val_in[1:0], f0val_in[1:0]}),
		.dout({error_stall, f2val[1:0], f1val[1:0], f0val[1:0]})
	);
	generate
		if (pt[2130-:5] == 1) begin
			rvdffe #(.WIDTH(BRDATA_SIZE)) brdata2ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[2]),
				.din(brdata_in[BRDATA_SIZE - 1:0]),
				.dout(brdata2[BRDATA_SIZE - 1:0])
			);
			rvdffe #(.WIDTH(BRDATA_SIZE)) brdata1ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[1]),
				.din(brdata_in[BRDATA_SIZE - 1:0]),
				.dout(brdata1[BRDATA_SIZE - 1:0])
			);
			rvdffe #(.WIDTH(BRDATA_SIZE)) brdata0ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[0]),
				.din(brdata_in[BRDATA_SIZE - 1:0]),
				.dout(brdata0[BRDATA_SIZE - 1:0])
			);
			rvdffe #(.WIDTH(MSIZE)) misc2ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[2]),
				.din(misc_data_in[MHI:0]),
				.dout(misc2[MHI:0])
			);
			rvdffe #(.WIDTH(MSIZE)) misc1ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[1]),
				.din(misc_data_in[MHI:0]),
				.dout(misc1[MHI:0])
			);
			rvdffe #(.WIDTH(MSIZE)) misc0ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(qwen[0]),
				.din(misc_data_in[MHI:0]),
				.dout(misc0[MHI:0])
			);
		end
		else rvdffie #(.WIDTH((MSIZE * 3) + (BRDATA_SIZE * 3))) miscff(
			.clk(clk),
			.rst_l(rst_l),
			.scan_mode(scan_mode),
			.din({(qwen[2] ? {misc_data_in[MHI:0], brdata_in[BRDATA_SIZE - 1:0]} : {misc2[MHI:0], brdata2[BRDATA_SIZE - 1:0]}), (qwen[1] ? {misc_data_in[MHI:0], brdata_in[BRDATA_SIZE - 1:0]} : {misc1[MHI:0], brdata1[BRDATA_SIZE - 1:0]}), (qwen[0] ? {misc_data_in[MHI:0], brdata_in[BRDATA_SIZE - 1:0]} : {misc0[MHI:0], brdata0[BRDATA_SIZE - 1:0]})}),
			.dout({misc2[MHI:0], misc1[MHI:0], misc0[MHI:0], brdata2[BRDATA_SIZE - 1:0], brdata1[BRDATA_SIZE - 1:0], brdata0[BRDATA_SIZE - 1:0]})
		);
	endgenerate
	wire [31:1] q2pc;
	wire [31:1] q1pc;
	wire [31:1] q0pc;
	rvdffe #(.WIDTH(31)) q2pcff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[2]),
		.din(ifu_fetch_pc[31:1]),
		.dout(q2pc[31:1])
	);
	rvdffe #(.WIDTH(31)) q1pcff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[1]),
		.din(ifu_fetch_pc[31:1]),
		.dout(q1pc[31:1])
	);
	rvdffe #(.WIDTH(31)) q0pcff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[0]),
		.din(ifu_fetch_pc[31:1]),
		.dout(q0pc[31:1])
	);
	rvdffe #(.WIDTH(32)) q2ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[2]),
		.din(ifu_fetch_data_f[31:0]),
		.dout(q2[31:0])
	);
	rvdffe #(.WIDTH(32)) q1ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[1]),
		.din(ifu_fetch_data_f[31:0]),
		.dout(q1[31:0])
	);
	rvdffe #(.WIDTH(32)) q0ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.en(qwen[0]),
		.din(ifu_fetch_data_f[31:0]),
		.dout(q0[31:0])
	);
	assign qren[2:0] = {rdptr[1:0] == 2'b10, rdptr[1:0] == 2'b01, rdptr[1:0] == 2'b00};
	assign qwen[2:0] = {(wrptr[1:0] == 2'b10) & ifvalid, (wrptr[1:0] == 2'b01) & ifvalid, (wrptr[1:0] == 2'b00) & ifvalid};
	assign rdptr_in[1:0] = (((((({2 {(qren[0] & ifu_fb_consume1) & ~exu_flush_final}} & 2'b01) | ({2 {(qren[1] & ifu_fb_consume1) & ~exu_flush_final}} & 2'b10)) | ({2 {(qren[2] & ifu_fb_consume1) & ~exu_flush_final}} & 2'b00)) | ({2 {(qren[0] & ifu_fb_consume2) & ~exu_flush_final}} & 2'b10)) | ({2 {(qren[1] & ifu_fb_consume2) & ~exu_flush_final}} & 2'b00)) | ({2 {(qren[2] & ifu_fb_consume2) & ~exu_flush_final}} & 2'b01)) | ({2 {(~ifu_fb_consume1 & ~ifu_fb_consume2) & ~exu_flush_final}} & rdptr[1:0]);
	assign wrptr_in[1:0] = ((({2 {qwen[0] & ~exu_flush_final}} & 2'b01) | ({2 {qwen[1] & ~exu_flush_final}} & 2'b10)) | ({2 {qwen[2] & ~exu_flush_final}} & 2'b00)) | ({2 {~ifvalid & ~exu_flush_final}} & wrptr[1:0]);
	assign q2off_in = (((~qwen[2] & (rdptr[1:0] == 2'd2)) & (q2off | f0_shift_2B)) | ((~qwen[2] & (rdptr[1:0] == 2'd1)) & (q2off | f1_shift_2B))) | ((~qwen[2] & (rdptr[1:0] == 2'd0)) & q2off);
	assign q1off_in = (((~qwen[1] & (rdptr[1:0] == 2'd1)) & (q1off | f0_shift_2B)) | ((~qwen[1] & (rdptr[1:0] == 2'd0)) & (q1off | f1_shift_2B))) | ((~qwen[1] & (rdptr[1:0] == 2'd2)) & q1off);
	assign q0off_in = (((~qwen[0] & (rdptr[1:0] == 2'd0)) & (q0off | f0_shift_2B)) | ((~qwen[0] & (rdptr[1:0] == 2'd2)) & (q0off | f1_shift_2B))) | ((~qwen[0] & (rdptr[1:0] == 2'd1)) & q0off);
	assign q0ptr = (((rdptr[1:0] == 2'b00) & q0off) | ((rdptr[1:0] == 2'b01) & q1off)) | ((rdptr[1:0] == 2'b10) & q2off);
	assign q1ptr = (((rdptr[1:0] == 2'b00) & q1off) | ((rdptr[1:0] == 2'b01) & q2off)) | ((rdptr[1:0] == 2'b10) & q0off);
	assign q0sel[1:0] = {q0ptr, ~q0ptr};
	assign q1sel[1:0] = {q1ptr, ~q1ptr};
	generate
		if (pt[2130-:5] == 1) begin
			assign misc_data_in[MHI:0] = {ic_access_fault_type_f[1:0], ifu_bp_btb_target_f[31:1], ifu_bp_poffset_f[11:0], ifu_bp_fghr_f[pt[2236-:8] - 1:0]};
		end
		else assign misc_data_in[MHI:0] = {ic_access_fault_type_f[1:0]};
	endgenerate
	assign {misc1eff[MHI:0], misc0eff[MHI:0]} = (({MSIZE * 2 {qren[0]}} & {misc1[MHI:0], misc0[MHI:0]}) | ({MSIZE * 2 {qren[1]}} & {misc2[MHI:0], misc1[MHI:0]})) | ({MSIZE * 2 {qren[2]}} & {misc0[MHI:0], misc2[MHI:0]});
	generate
		if (pt[2130-:5] == 1) begin
			assign {f1ictype[1:0], f1prett[31:1], f1poffset[11:0], f1fghr[pt[2236-:8] - 1:0]} = misc1eff[MHI:0];
			assign {f0ictype[1:0], f0prett[31:1], f0poffset[11:0], f0fghr[pt[2236-:8] - 1:0]} = misc0eff[MHI:0];
			if (pt[2120-:5]) begin
				assign brdata_in[BRDATA_SIZE - 1:0] = {ifu_bp_fa_index_f[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])], iccm_rd_ecc_double_err[1], ic_access_fault_f[1], ifu_bp_hist1_f[1], ifu_bp_hist0_f[1], ifu_bp_pc4_f[1], ifu_bp_way_f[1], ifu_bp_valid_f[1], ifu_bp_ret_f[1], ifu_bp_fa_index_f[0+:$clog2(pt[2061-:14])], iccm_rd_ecc_double_err[0], ic_access_fault_f[0], ifu_bp_hist1_f[0], ifu_bp_hist0_f[0], ifu_bp_pc4_f[0], ifu_bp_way_f[0], ifu_bp_valid_f[0], ifu_bp_ret_f[0]};
				assign {f0index[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])], f0dbecc[1], f0icaf[1], f0hist1[1], f0hist0[1], f0pc4[1], f0way[1], f0brend[1], f0ret[1], f0index[0+:$clog2(pt[2061-:14])], f0dbecc[0], f0icaf[0], f0hist1[0], f0hist0[0], f0pc4[0], f0way[0], f0brend[0], f0ret[0]} = brdata0final[BRDATA_SIZE - 1:0];
				assign {f1index[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])], f1dbecc[1], f1icaf[1], f1hist1[1], f1hist0[1], f1pc4[1], f1way[1], f1brend[1], f1ret[1], f1index[0+:$clog2(pt[2061-:14])], f1dbecc[0], f1icaf[0], f1hist1[0], f1hist0[0], f1pc4[0], f1way[0], f1brend[0], f1ret[0]} = brdata1final[BRDATA_SIZE - 1:0];
			end
			else begin
				assign brdata_in[BRDATA_SIZE - 1:0] = {iccm_rd_ecc_double_err[1], ic_access_fault_f[1], ifu_bp_hist1_f[1], ifu_bp_hist0_f[1], ifu_bp_pc4_f[1], ifu_bp_way_f[1], ifu_bp_valid_f[1], ifu_bp_ret_f[1], iccm_rd_ecc_double_err[0], ic_access_fault_f[0], ifu_bp_hist1_f[0], ifu_bp_hist0_f[0], ifu_bp_pc4_f[0], ifu_bp_way_f[0], ifu_bp_valid_f[0], ifu_bp_ret_f[0]};
				assign {f0dbecc[1], f0icaf[1], f0hist1[1], f0hist0[1], f0pc4[1], f0way[1], f0brend[1], f0ret[1], f0dbecc[0], f0icaf[0], f0hist1[0], f0hist0[0], f0pc4[0], f0way[0], f0brend[0], f0ret[0]} = brdata0final[BRDATA_SIZE - 1:0];
				assign {f1dbecc[1], f1icaf[1], f1hist1[1], f1hist0[1], f1pc4[1], f1way[1], f1brend[1], f1ret[1], f1dbecc[0], f1icaf[0], f1hist1[0], f1hist0[0], f1pc4[0], f1way[0], f1brend[0], f1ret[0]} = brdata1final[BRDATA_SIZE - 1:0];
			end
			assign {brdata1eff[BRDATA_SIZE - 1:0], brdata0eff[BRDATA_SIZE - 1:0]} = (({BRDATA_SIZE * 2 {qren[0]}} & {brdata1[BRDATA_SIZE - 1:0], brdata0[BRDATA_SIZE - 1:0]}) | ({BRDATA_SIZE * 2 {qren[1]}} & {brdata2[BRDATA_SIZE - 1:0], brdata1[BRDATA_SIZE - 1:0]})) | ({BRDATA_SIZE * 2 {qren[2]}} & {brdata0[BRDATA_SIZE - 1:0], brdata2[BRDATA_SIZE - 1:0]});
			assign brdata0final[BRDATA_SIZE - 1:0] = ({BRDATA_SIZE {q0sel[0]}} & {brdata0eff[(2 * BRDATA_WIDTH) - 1:0]}) | ({BRDATA_SIZE {q0sel[1]}} & {{BRDATA_WIDTH {1'b0}}, brdata0eff[BRDATA_SIZE - 1:BRDATA_WIDTH]});
			assign brdata1final[BRDATA_SIZE - 1:0] = ({BRDATA_SIZE {q1sel[0]}} & {brdata1eff[(2 * BRDATA_WIDTH) - 1:0]}) | ({BRDATA_SIZE {q1sel[1]}} & {{BRDATA_WIDTH {1'b0}}, brdata1eff[BRDATA_SIZE - 1:BRDATA_WIDTH]});
		end
		else begin
			assign {f1ictype[1:0]} = misc1eff[MHI:0];
			assign {f0ictype[1:0]} = misc0eff[MHI:0];
			assign brdata_in[BRDATA_SIZE - 1:0] = {iccm_rd_ecc_double_err[1], ic_access_fault_f[1], iccm_rd_ecc_double_err[0], ic_access_fault_f[0]};
			assign {f0dbecc[1], f0icaf[1], f0dbecc[0], f0icaf[0]} = brdata0final[BRDATA_SIZE - 1:0];
			assign {f1dbecc[1], f1icaf[1], f1dbecc[0], f1icaf[0]} = brdata1final[BRDATA_SIZE - 1:0];
			assign {brdata1eff[BRDATA_SIZE - 1:0], brdata0eff[BRDATA_SIZE - 1:0]} = (({BRDATA_SIZE * 2 {qren[0]}} & {brdata1[BRDATA_SIZE - 1:0], brdata0[BRDATA_SIZE - 1:0]}) | ({BRDATA_SIZE * 2 {qren[1]}} & {brdata2[BRDATA_SIZE - 1:0], brdata1[BRDATA_SIZE - 1:0]})) | ({BRDATA_SIZE * 2 {qren[2]}} & {brdata0[BRDATA_SIZE - 1:0], brdata2[BRDATA_SIZE - 1:0]});
			assign brdata0final[BRDATA_SIZE - 1:0] = ({BRDATA_SIZE {q0sel[0]}} & {brdata0eff[(2 * BRDATA_WIDTH) - 1:0]}) | ({BRDATA_SIZE {q0sel[1]}} & {{BRDATA_WIDTH {1'b0}}, brdata0eff[BRDATA_SIZE - 1:BRDATA_WIDTH]});
			assign brdata1final[BRDATA_SIZE - 1:0] = ({BRDATA_SIZE {q1sel[0]}} & {brdata1eff[(2 * BRDATA_WIDTH) - 1:0]}) | ({BRDATA_SIZE {q1sel[1]}} & {{BRDATA_WIDTH {1'b0}}, brdata1eff[BRDATA_SIZE - 1:BRDATA_WIDTH]});
		end
	endgenerate
	assign f2_valid = f2val[0];
	assign sf1_valid = sf1val[0];
	assign sf0_valid = sf0val[0];
	assign consume_fb0 = ~sf0val[0] & f0val[0];
	assign consume_fb1 = ~sf1val[0] & f1val[0];
	assign ifu_fb_consume1 = (consume_fb0 & ~consume_fb1) & ~exu_flush_final;
	assign ifu_fb_consume2 = (consume_fb0 & consume_fb1) & ~exu_flush_final;
	assign ifvalid = ifu_fetch_val[0];
	assign shift_f1_f0 = ~sf0_valid & sf1_valid;
	assign shift_f2_f0 = (~sf0_valid & ~sf1_valid) & f2_valid;
	assign shift_f2_f1 = (~sf0_valid & sf1_valid) & f2_valid;
	assign fetch_to_f0 = ((~sf0_valid & ~sf1_valid) & ~f2_valid) & ifvalid;
	assign fetch_to_f1 = ((((~sf0_valid & ~sf1_valid) & f2_valid) & ifvalid) | (((~sf0_valid & sf1_valid) & ~f2_valid) & ifvalid)) | (((sf0_valid & ~sf1_valid) & ~f2_valid) & ifvalid);
	assign fetch_to_f2 = (((~sf0_valid & sf1_valid) & f2_valid) & ifvalid) | (((sf0_valid & sf1_valid) & ~f2_valid) & ifvalid);
	assign f2val_in[1:0] = ({2 {fetch_to_f2 & ~exu_flush_final}} & ifu_fetch_val[1:0]) | ({2 {((~fetch_to_f2 & ~shift_f2_f1) & ~shift_f2_f0) & ~exu_flush_final}} & f2val[1:0]);
	assign sf1val[1:0] = ({2 {f1_shift_2B}} & {1'b0, f1val[1]}) | ({2 {~f1_shift_2B}} & f1val[1:0]);
	assign f1val_in[1:0] = (({2 {fetch_to_f1 & ~exu_flush_final}} & ifu_fetch_val[1:0]) | ({2 {shift_f2_f1 & ~exu_flush_final}} & f2val[1:0])) | ({2 {((~fetch_to_f1 & ~shift_f2_f1) & ~shift_f1_f0) & ~exu_flush_final}} & sf1val[1:0]);
	assign sf0val[1:0] = ({2 {shift_2B}} & {1'b0, f0val[1]}) | ({2 {~shift_2B & ~shift_4B}} & f0val[1:0]);
	assign f0val_in[1:0] = ((({2 {fetch_to_f0 & ~exu_flush_final}} & ifu_fetch_val[1:0]) | ({2 {shift_f2_f0 & ~exu_flush_final}} & f2val[1:0])) | ({2 {shift_f1_f0 & ~exu_flush_final}} & sf1val[1:0])) | ({2 {((~fetch_to_f0 & ~shift_f2_f0) & ~shift_f1_f0) & ~exu_flush_final}} & sf0val[1:0]);
	assign {q1eff[31:0], q0eff[31:0]} = (({64 {qren[0]}} & {q1[31:0], q0[31:0]}) | ({64 {qren[1]}} & {q2[31:0], q1[31:0]})) | ({64 {qren[2]}} & {q0[31:0], q2[31:0]});
	assign q0final[31:0] = ({32 {q0sel[0]}} & {q0eff[31:0]}) | ({32 {q0sel[1]}} & {16'b0000000000000000, q0eff[31:16]});
	assign q1final[15:0] = ({16 {q1sel[0]}} & q1eff[15:0]) | ({16 {q1sel[1]}} & q1eff[31:16]);
	wire [31:1] q0pceff;
	wire [31:1] q0pcfinal;
	wire [31:1] q1pceff;
	assign {q1pceff[31:1], q0pceff[31:1]} = (({62 {qren[0]}} & {q1pc[31:1], q0pc[31:1]}) | ({62 {qren[1]}} & {q2pc[31:1], q1pc[31:1]})) | ({62 {qren[2]}} & {q0pc[31:1], q2pc[31:1]});
	assign q0pcfinal[31:1] = ({31 {q0sel[0]}} & q0pceff[31:1]) | ({31 {q0sel[1]}} & (q0pceff[31:1] + 31'd1));
	assign aligndata[31:0] = ({32 {f0val[1]}} & {q0final[31:0]}) | ({32 {~f0val[1] & f0val[0]}} & {q1final[15:0], q0final[15:0]});
	assign alignval[1:0] = ({2 {f0val[1]}} & 2'b11) | ({2 {~f0val[1] & f0val[0]}} & {f1val[0], 1'b1});
	assign alignicaf[1:0] = ({2 {f0val[1]}} & f0icaf[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1icaf[0], f0icaf[0]});
	assign aligndbecc[1:0] = ({2 {f0val[1]}} & f0dbecc[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1dbecc[0], f0dbecc[0]});
	generate
		if (pt[2130-:5] == 1) begin
			assign alignbrend[1:0] = ({2 {f0val[1]}} & f0brend[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1brend[0], f0brend[0]});
			assign alignpc4[1:0] = ({2 {f0val[1]}} & f0pc4[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1pc4[0], f0pc4[0]});
			if (pt[2120-:5]) begin
				assign alignindex[0+:$clog2(pt[2061-:14])] = f0index[0+:$clog2(pt[2061-:14])];
				assign alignindex[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])] = (f0val[1] ? f0index[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])] : f1index[0+:$clog2(pt[2061-:14])]);
			end
			assign alignret[1:0] = ({2 {f0val[1]}} & f0ret[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1ret[0], f0ret[0]});
			assign alignway[1:0] = ({2 {f0val[1]}} & f0way[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1way[0], f0way[0]});
			assign alignhist1[1:0] = ({2 {f0val[1]}} & f0hist1[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1hist1[0], f0hist1[0]});
			assign alignhist0[1:0] = ({2 {f0val[1]}} & f0hist0[1:0]) | ({2 {~f0val[1] & f0val[0]}} & {f1hist0[0], f0hist0[0]});
			assign secondpc[31:1] = ({31 {f0val[1]}} & (q0pceff[31:1] + 31'd1)) | ({31 {~f0val[1] & f0val[0]}} & q1pceff[31:1]);
			assign firstpc[31:1] = q0pcfinal[31:1];
		end
	endgenerate
	assign alignfromf1[1] = ~f0val[1] & f0val[0];
	assign ifu_i0_pc[31:1] = q0pcfinal[31:1];
	assign ifu_i0_pc4 = first4B;
	assign ifu_i0_cinst[15:0] = aligndata[15:0];
	assign first4B = aligndata[1:0] == 2'b11;
	assign first2B = ~first4B;
	assign ifu_i0_valid = (first4B & alignval[1]) | (first2B & alignval[0]);
	assign ifu_i0_icaf = (first4B & |alignicaf[1:0]) | (first2B & alignicaf[0]);
	assign ifu_i0_icaf_type[1:0] = ((((first4B & ~f0val[1]) & f0val[0]) & ~alignicaf[0]) & ~aligndbecc[0] ? f1ictype[1:0] : f0ictype[1:0]);
	assign icaf_eff[1:0] = alignicaf[1:0] | aligndbecc[1:0];
	assign ifu_i0_icaf_second = (first4B & ~icaf_eff[0]) & icaf_eff[1];
	assign ifu_i0_dbecc = (first4B & |aligndbecc[1:0]) | (first2B & aligndbecc[0]);
	assign ifirst[31:0] = aligndata[31:0];
	assign ifu_i0_instr[31:0] = ({32 {first4B & alignval[1]}} & ifirst[31:0]) | ({32 {first2B & alignval[0]}} & uncompress0[31:0]);
	generate
		if (pt[2130-:5] == 1) begin
			eb1_btb_addr_hash #(.pt(pt)) firsthash(
				.pc(firstpc[pt[2079-:9]:pt[2106-:9]]),
				.hash(firstpc_hash[pt[2172-:9]:pt[2163-:6]])
			);
			eb1_btb_addr_hash #(.pt(pt)) secondhash(
				.pc(secondpc[pt[2079-:9]:pt[2106-:9]]),
				.hash(secondpc_hash[pt[2172-:9]:pt[2163-:6]])
			);
			if (pt[2120-:5]) begin
				assign firstbrtag_hash = firstpc;
				assign secondbrtag_hash = secondpc;
			end
			else if (pt[2144-:5]) begin : btbfold
				eb1_btb_tag_hash_fold #(.pt(pt)) first_brhash(
					.pc(firstpc[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]),
					.hash(firstbrtag_hash[pt[2139-:9] - 1:0])
				);
				eb1_btb_tag_hash_fold #(.pt(pt)) second_brhash(
					.pc(secondpc[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]),
					.hash(secondbrtag_hash[pt[2139-:9] - 1:0])
				);
			end
			else begin
				eb1_btb_tag_hash #(.pt(pt)) first_brhash(
					.pc(firstpc[((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]),
					.hash(firstbrtag_hash[pt[2139-:9] - 1:0])
				);
				eb1_btb_tag_hash #(.pt(pt)) second_brhash(
					.pc(secondpc[((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]),
					.hash(secondbrtag_hash[pt[2139-:9] - 1:0])
				);
			end
			always @(*) begin
				i0_brp = {51 {1'sb0}};
				i0_br_start_error = (first4B & alignval[1]) & alignbrend[0];
				i0_brp[50] = ((first2B & alignbrend[0]) | (first4B & alignbrend[1])) | i0_br_start_error;
				i0_brp_pc4 = (first2B & alignpc4[0]) | (first4B & alignpc4[1]);
				i0_brp[0] = (first2B & alignret[0]) | (first4B & alignret[1]);
				i0_brp[1] = (first2B | alignbrend[0] ? alignway[0] : alignway[1]);
				i0_brp[37] = (first2B & alignhist1[0]) | (first4B & alignhist1[1]);
				i0_brp[36] = (first2B & alignhist0[0]) | (first4B & alignhist0[1]);
				i0_ends_f1 = first4B & alignfromf1[1];
				i0_brp[49:38] = (i0_ends_f1 ? f1poffset[11:0] : f0poffset[11:0]);
				i0_brp[32:2] = (i0_ends_f1 ? f1prett[31:1] : f0prett[31:1]);
				i0_brp[34] = i0_br_start_error;
				i0_brp[33] = (first2B | alignbrend[0] ? firstpc[1] : secondpc[1]);
				i0_brp[35] = ((i0_brp[50] & i0_brp_pc4) & first2B) | ((i0_brp[50] & ~i0_brp_pc4) & first4B);
				if (pt[2120-:5])
					ifu_i0_fa_index = (first2B | alignbrend[0] ? alignindex[0+:$clog2(pt[2061-:14])] : alignindex[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])]);
				else
					ifu_i0_fa_index = {$clog2(pt[2061-:14]) {1'sb0}};
			end
			assign ifu_i0_bp_index[pt[2172-:9]:pt[2163-:6]] = (first2B | alignbrend[0] ? firstpc_hash[pt[2172-:9]:pt[2163-:6]] : secondpc_hash[pt[2172-:9]:pt[2163-:6]]);
			assign ifu_i0_bp_fghr[pt[2236-:8] - 1:0] = (i0_ends_f1 ? f1fghr[pt[2236-:8] - 1:0] : f0fghr[pt[2236-:8] - 1:0]);
			assign ifu_i0_bp_btag[pt[2139-:9] - 1:0] = (first2B | alignbrend[0] ? firstbrtag_hash[pt[2139-:9] - 1:0] : secondbrtag_hash[pt[2139-:9] - 1:0]);
		end
		else begin
			wire [51:1] sv2v_tmp_B43E9;
			assign sv2v_tmp_B43E9 = {51 {1'sb0}};
			always @(*) i0_brp = sv2v_tmp_B43E9;
			assign ifu_i0_bp_index = {(pt[2172-:9] >= pt[2163-:6] ? (pt[2172-:9] - pt[2163-:6]) + 1 : (pt[2163-:6] - pt[2172-:9]) + 1) {1'sb0}};
			assign ifu_i0_bp_fghr = {pt[2236-:8] {1'sb0}};
			assign ifu_i0_bp_btag = {pt[2139-:9] {1'sb0}};
		end
	endgenerate
	eb1_ifu_compress_ctl #(.pt(pt)) compress0(
		.din((first2B ? aligndata[15:0] : {16 {1'sb0}})),
		.dout(uncompress0[31:0])
	);
	assign i0_shift = dec_i0_decode_d & ~error_stall;
	assign ifu_pmu_instr_aligned = i0_shift;
	assign shift_2B = i0_shift & first2B;
	assign shift_4B = i0_shift & first4B;
	assign f0_shift_2B = (shift_2B & f0val[0]) | ((shift_4B & f0val[0]) & ~f0val[1]);
	assign f1_shift_2B = (f0val[0] & ~f0val[1]) & shift_4B;
endmodule
module eb1_ifu_bp_ctl (
	clk,
	rst_l,
	ic_hit_f,
	ifc_fetch_addr_f,
	ifc_fetch_req_f,
	dec_tlu_br0_r_pkt,
	exu_i0_br_fghr_r,
	exu_i0_br_index_r,
	dec_fa_error_index,
	dec_tlu_flush_lower_wb,
	dec_tlu_flush_leak_one_wb,
	dec_tlu_bpred_disable,
	exu_mp_pkt,
	exu_mp_eghr,
	exu_mp_fghr,
	exu_mp_index,
	exu_mp_btag,
	exu_flush_final,
	ifu_bp_hit_taken_f,
	ifu_bp_btb_target_f,
	ifu_bp_inst_mask_f,
	ifu_bp_fghr_f,
	ifu_bp_way_f,
	ifu_bp_ret_f,
	ifu_bp_hist1_f,
	ifu_bp_hist0_f,
	ifu_bp_pc4_f,
	ifu_bp_valid_f,
	ifu_bp_poffset_f,
	ifu_bp_fa_index_f,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire ic_hit_f;
	input wire [31:1] ifc_fetch_addr_f;
	input wire ifc_fetch_req_f;
	input wire [6:0] dec_tlu_br0_r_pkt;
	input wire [pt[2236-:8] - 1:0] exu_i0_br_fghr_r;
	input wire [pt[2172-:9]:pt[2163-:6]] exu_i0_br_index_r;
	input wire [$clog2(pt[2061-:14]) - 1:0] dec_fa_error_index;
	input wire dec_tlu_flush_lower_wb;
	input wire dec_tlu_flush_leak_one_wb;
	input wire dec_tlu_bpred_disable;
	input wire [55:0] exu_mp_pkt;
	input wire [pt[2236-:8] - 1:0] exu_mp_eghr;
	input wire [pt[2236-:8] - 1:0] exu_mp_fghr;
	input wire [pt[2172-:9]:pt[2163-:6]] exu_mp_index;
	input wire [pt[2139-:9] - 1:0] exu_mp_btag;
	input wire exu_flush_final;
	output wire ifu_bp_hit_taken_f;
	output wire [31:1] ifu_bp_btb_target_f;
	output wire ifu_bp_inst_mask_f;
	output wire [pt[2236-:8] - 1:0] ifu_bp_fghr_f;
	output wire [1:0] ifu_bp_way_f;
	output wire [1:0] ifu_bp_ret_f;
	output wire [1:0] ifu_bp_hist1_f;
	output wire [1:0] ifu_bp_hist0_f;
	output wire [1:0] ifu_bp_pc4_f;
	output wire [1:0] ifu_bp_valid_f;
	output wire [11:0] ifu_bp_poffset_f;
	output wire [(2 * $clog2(pt[2061-:14])) - 1:0] ifu_bp_fa_index_f;
	input wire scan_mode;
	localparam BTB_DWIDTH = (pt[2047-:9] + pt[2139-:9]) + 5;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	localparam BTB_DWIDTH_TOP = (sv2v_cast_32_signed(pt[2047-:9]) + sv2v_cast_32_signed(pt[2139-:9])) + 4;
	localparam BTB_FA_INDEX = $clog2(pt[2061-:14]) - 1;
	localparam FA_CMP_LOWER = $clog2(pt[1095-:11]);
	localparam FA_TAG_END_UPPER = ((5 + sv2v_cast_32_signed(pt[2047-:9])) + FA_CMP_LOWER) - 1;
	localparam FA_TAG_START_LOWER = (3 + sv2v_cast_32_signed(pt[2047-:9])) + FA_CMP_LOWER;
	localparam FA_TAG_END_LOWER = 5 + sv2v_cast_32_signed(pt[2047-:9]);
	localparam TAG_START = BTB_DWIDTH - 1;
	localparam PC4 = 4;
	localparam BOFF = 3;
	localparam CALL = 2;
	localparam RET = 1;
	localparam BV = 0;
	localparam LRU_SIZE = pt[2157-:13];
	localparam NUM_BHT_LOOP = (pt[2256-:15] > 16 ? 16 : pt[2256-:15]);
	localparam NUM_BHT_LOOP_INNER_HI = (pt[2256-:15] > 16 ? pt[2262-:6] + 3 : pt[2270-:8]);
	localparam NUM_BHT_LOOP_OUTER_LO = (pt[2256-:15] > 16 ? pt[2262-:6] + 4 : pt[2262-:6]);
	localparam BHT_NO_ADDR_MATCH = pt[2256-:15] <= 16;
	wire exu_mp_valid_write;
	wire exu_mp_ataken;
	wire exu_mp_valid;
	wire exu_mp_boffset;
	wire exu_mp_pc4;
	wire exu_mp_call;
	wire exu_mp_ret;
	wire exu_mp_ja;
	wire [1:0] exu_mp_hist;
	wire [11:0] exu_mp_tgt;
	wire [pt[2172-:9]:pt[2163-:6]] exu_mp_addr;
	wire dec_tlu_br0_v_wb;
	wire [1:0] dec_tlu_br0_hist_wb;
	wire [pt[2172-:9]:pt[2163-:6]] dec_tlu_br0_addr_wb;
	wire dec_tlu_br0_error_wb;
	wire dec_tlu_br0_start_error_wb;
	wire [pt[2236-:8] - 1:0] exu_i0_br_fghr_wb;
	wire use_mp_way;
	wire use_mp_way_p1;
	wire [(pt[31-:8] * 32) - 1:0] rets_out;
	wire [(pt[31-:8] * 32) - 1:0] rets_in;
	wire [pt[31-:8] - 1:0] rsenable;
	wire [11:0] btb_rd_tgt_f;
	wire btb_rd_pc4_f;
	wire btb_rd_call_f;
	wire btb_rd_ret_f;
	wire [1:1] bp_total_branch_offset_f;
	wire [31:1] bp_btb_target_adder_f;
	wire [31:1] bp_rs_call_target_f;
	wire rs_push;
	wire rs_pop;
	wire rs_hold;
	wire [pt[2172-:9]:pt[2163-:6]] btb_rd_addr_p1_f;
	wire [pt[2172-:9]:pt[2163-:6]] btb_wr_addr;
	wire [pt[2172-:9]:pt[2163-:6]] btb_rd_addr_f;
	wire [pt[2139-:9] - 1:0] btb_wr_tag;
	wire [pt[2139-:9] - 1:0] fetch_rd_tag_f;
	wire [pt[2139-:9] - 1:0] fetch_rd_tag_p1_f;
	wire [BTB_DWIDTH - 1:0] btb_wr_data;
	wire btb_wr_en_way0;
	wire btb_wr_en_way1;
	wire dec_tlu_error_wb;
	wire btb_valid;
	wire dec_tlu_br0_middle_wb;
	wire [pt[2172-:9]:pt[2163-:6]] btb_error_addr_wb;
	wire branch_error_collision_f;
	wire fetch_mp_collision_f;
	wire branch_error_collision_p1_f;
	wire fetch_mp_collision_p1_f;
	wire branch_error_bank_conflict_f;
	wire [pt[2236-:8] - 1:0] merged_ghr;
	wire [pt[2236-:8] - 1:0] fghr_ns;
	wire [pt[2236-:8] - 1:0] fghr;
	wire [1:0] num_valids;
	wire [LRU_SIZE - 1:0] btb_lru_b0_f;
	wire [LRU_SIZE - 1:0] btb_lru_b0_hold;
	wire [LRU_SIZE - 1:0] btb_lru_b0_ns;
	wire [LRU_SIZE - 1:0] fetch_wrindex_dec;
	wire [LRU_SIZE - 1:0] fetch_wrindex_p1_dec;
	wire [LRU_SIZE - 1:0] fetch_wrlru_b0;
	wire [LRU_SIZE - 1:0] fetch_wrlru_p1_b0;
	wire [LRU_SIZE - 1:0] mp_wrindex_dec;
	wire [LRU_SIZE - 1:0] mp_wrlru_b0;
	wire btb_lru_rd_f;
	wire btb_lru_rd_p1_f;
	wire lru_update_valid_f;
	wire tag_match_way0_f;
	wire tag_match_way1_f;
	wire [1:0] way_raw;
	wire [1:0] bht_dir_f;
	wire [1:0] btb_sel_f;
	wire [1:0] wayhit_f;
	wire [1:0] vwayhit_f;
	wire [1:0] wayhit_p1_f;
	wire [1:0] bht_valid_f;
	wire [1:0] bht_force_taken_f;
	wire leak_one_f;
	wire leak_one_f_d1;
	wire [(LRU_SIZE * BTB_DWIDTH) - 1:0] btb_bank0_rd_data_way0_out;
	wire [(LRU_SIZE * BTB_DWIDTH) - 1:0] btb_bank0_rd_data_way1_out;
	reg [BTB_DWIDTH - 1:0] btb_bank0_rd_data_way0_f;
	reg [BTB_DWIDTH - 1:0] btb_bank0_rd_data_way1_f;
	reg [BTB_DWIDTH - 1:0] btb_bank0_rd_data_way0_p1_f;
	reg [BTB_DWIDTH - 1:0] btb_bank0_rd_data_way1_p1_f;
	reg [BTB_DWIDTH - 1:0] btb_vbank0_rd_data_f;
	reg [BTB_DWIDTH - 1:0] btb_vbank1_rd_data_f;
	wire final_h;
	wire btb_fg_crossing_f;
	wire middle_of_bank;
	wire [1:0] bht_vbank0_rd_data_f;
	wire [1:0] bht_vbank1_rd_data_f;
	wire branch_error_bank_conflict_p1_f;
	wire tag_match_way0_p1_f;
	wire tag_match_way1_p1_f;
	wire [1:0] btb_vlru_rd_f;
	wire [1:0] fetch_start_f;
	wire [1:0] tag_match_vway1_expanded_f;
	wire [1:0] tag_match_way0_expanded_p1_f;
	wire [1:0] tag_match_way1_expanded_p1_f;
	wire [31:2] fetch_addr_p1_f;
	wire exu_mp_way;
	wire exu_mp_way_f;
	wire dec_tlu_br0_way_wb;
	wire dec_tlu_way_wb;
	wire [BTB_DWIDTH - 1:0] btb_bank0e_rd_data_f;
	wire [BTB_DWIDTH - 1:0] btb_bank0e_rd_data_p1_f;
	wire [BTB_DWIDTH - 1:0] btb_bank0o_rd_data_f;
	wire [1:0] tag_match_way0_expanded_f;
	wire [1:0] tag_match_way1_expanded_f;
	reg [1:0] bht_bank0_rd_data_f;
	reg [1:0] bht_bank1_rd_data_f;
	reg [1:0] bht_bank0_rd_data_p1_f;
	genvar j;
	genvar i;
	assign exu_mp_valid = exu_mp_pkt[55] & ~leak_one_f;
	assign exu_mp_boffset = exu_mp_pkt[53];
	assign exu_mp_pc4 = exu_mp_pkt[52];
	assign exu_mp_call = exu_mp_pkt[34];
	assign exu_mp_ret = exu_mp_pkt[31];
	assign exu_mp_ja = exu_mp_pkt[33];
	assign exu_mp_way = exu_mp_pkt[32];
	assign exu_mp_hist[1:0] = exu_mp_pkt[51:50];
	assign exu_mp_tgt[11:0] = exu_mp_pkt[49:38];
	assign exu_mp_addr[pt[2172-:9]:pt[2163-:6]] = exu_mp_index[pt[2172-:9]:pt[2163-:6]];
	assign exu_mp_ataken = exu_mp_pkt[54];
	assign dec_tlu_br0_v_wb = dec_tlu_br0_r_pkt[6];
	assign dec_tlu_br0_hist_wb[1:0] = dec_tlu_br0_r_pkt[5:4];
	assign dec_tlu_br0_addr_wb[pt[2172-:9]:pt[2163-:6]] = exu_i0_br_index_r[pt[2172-:9]:pt[2163-:6]];
	assign dec_tlu_br0_error_wb = dec_tlu_br0_r_pkt[3];
	assign dec_tlu_br0_middle_wb = dec_tlu_br0_r_pkt[0];
	assign dec_tlu_br0_way_wb = dec_tlu_br0_r_pkt[1];
	assign dec_tlu_br0_start_error_wb = dec_tlu_br0_r_pkt[2];
	assign exu_i0_br_fghr_wb[pt[2236-:8] - 1:0] = exu_i0_br_fghr_r[pt[2236-:8] - 1:0];
	eb1_btb_addr_hash #(.pt(pt)) f1hash(
		.pc(ifc_fetch_addr_f[pt[2079-:9]:pt[2106-:9]]),
		.hash(btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]])
	);
	assign fetch_addr_p1_f[31:2] = ifc_fetch_addr_f[31:2] + 30'b000000000000000000000000000001;
	eb1_btb_addr_hash #(.pt(pt)) f1hash_p1(
		.pc(fetch_addr_p1_f[pt[2079-:9]:pt[2106-:9]]),
		.hash(btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]])
	);
	assign btb_sel_f[1] = ~bht_dir_f[0];
	assign btb_sel_f[0] = bht_dir_f[0];
	assign fetch_start_f[1:0] = {ifc_fetch_addr_f[1], ~ifc_fetch_addr_f[1]};
	assign branch_error_collision_f = dec_tlu_error_wb & (btb_error_addr_wb[pt[2172-:9]:pt[2163-:6]] == btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]]);
	assign branch_error_collision_p1_f = dec_tlu_error_wb & (btb_error_addr_wb[pt[2172-:9]:pt[2163-:6]] == btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]]);
	assign branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb;
	assign branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb;
	assign leak_one_f = (dec_tlu_flush_leak_one_wb & dec_tlu_flush_lower_wb) | (leak_one_f_d1 & ~dec_tlu_flush_lower_wb);
	wire exu_flush_final_d1;
	generate
		if (!pt[2120-:5]) begin
			assign fetch_mp_collision_f = (((exu_mp_btag[pt[2139-:9] - 1:0] == fetch_rd_tag_f[pt[2139-:9] - 1:0]) & exu_mp_valid) & ifc_fetch_req_f) & (exu_mp_addr[pt[2172-:9]:pt[2163-:6]] == btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]]);
			assign fetch_mp_collision_p1_f = (((exu_mp_btag[pt[2139-:9] - 1:0] == fetch_rd_tag_p1_f[pt[2139-:9] - 1:0]) & exu_mp_valid) & ifc_fetch_req_f) & (exu_mp_addr[pt[2172-:9]:pt[2163-:6]] == btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]]);
			assign tag_match_way0_f = (((btb_bank0_rd_data_way0_f[BV] & (btb_bank0_rd_data_way0_f[TAG_START:17] == fetch_rd_tag_f[pt[2139-:9] - 1:0])) & ~(dec_tlu_way_wb & branch_error_bank_conflict_f)) & ifc_fetch_req_f) & ~leak_one_f;
			assign tag_match_way1_f = (((btb_bank0_rd_data_way1_f[BV] & (btb_bank0_rd_data_way1_f[TAG_START:17] == fetch_rd_tag_f[pt[2139-:9] - 1:0])) & ~(dec_tlu_way_wb & branch_error_bank_conflict_f)) & ifc_fetch_req_f) & ~leak_one_f;
			assign tag_match_way0_p1_f = (((btb_bank0_rd_data_way0_p1_f[BV] & (btb_bank0_rd_data_way0_p1_f[TAG_START:17] == fetch_rd_tag_p1_f[pt[2139-:9] - 1:0])) & ~(dec_tlu_way_wb & branch_error_bank_conflict_p1_f)) & ifc_fetch_req_f) & ~leak_one_f;
			assign tag_match_way1_p1_f = (((btb_bank0_rd_data_way1_p1_f[BV] & (btb_bank0_rd_data_way1_p1_f[TAG_START:17] == fetch_rd_tag_p1_f[pt[2139-:9] - 1:0])) & ~(dec_tlu_way_wb & branch_error_bank_conflict_p1_f)) & ifc_fetch_req_f) & ~leak_one_f;
			assign tag_match_way0_expanded_f[1:0] = {tag_match_way0_f & (btb_bank0_rd_data_way0_f[BOFF] ^ btb_bank0_rd_data_way0_f[PC4]), tag_match_way0_f & ~(btb_bank0_rd_data_way0_f[BOFF] ^ btb_bank0_rd_data_way0_f[PC4])};
			assign tag_match_way1_expanded_f[1:0] = {tag_match_way1_f & (btb_bank0_rd_data_way1_f[BOFF] ^ btb_bank0_rd_data_way1_f[PC4]), tag_match_way1_f & ~(btb_bank0_rd_data_way1_f[BOFF] ^ btb_bank0_rd_data_way1_f[PC4])};
			assign tag_match_way0_expanded_p1_f[1:0] = {tag_match_way0_p1_f & (btb_bank0_rd_data_way0_p1_f[BOFF] ^ btb_bank0_rd_data_way0_p1_f[PC4]), tag_match_way0_p1_f & ~(btb_bank0_rd_data_way0_p1_f[BOFF] ^ btb_bank0_rd_data_way0_p1_f[PC4])};
			assign tag_match_way1_expanded_p1_f[1:0] = {tag_match_way1_p1_f & (btb_bank0_rd_data_way1_p1_f[BOFF] ^ btb_bank0_rd_data_way1_p1_f[PC4]), tag_match_way1_p1_f & ~(btb_bank0_rd_data_way1_p1_f[BOFF] ^ btb_bank0_rd_data_way1_p1_f[PC4])};
			assign wayhit_f[1:0] = tag_match_way0_expanded_f[1:0] | tag_match_way1_expanded_f[1:0];
			assign wayhit_p1_f[1:0] = tag_match_way0_expanded_p1_f[1:0] | tag_match_way1_expanded_p1_f[1:0];
			assign btb_bank0o_rd_data_f[BTB_DWIDTH - 1:0] = ({17 + pt[2139-:9] {tag_match_way0_expanded_f[1]}} & btb_bank0_rd_data_way0_f[BTB_DWIDTH - 1:0]) | ({17 + pt[2139-:9] {tag_match_way1_expanded_f[1]}} & btb_bank0_rd_data_way1_f[BTB_DWIDTH - 1:0]);
			assign btb_bank0e_rd_data_f[BTB_DWIDTH - 1:0] = ({17 + pt[2139-:9] {tag_match_way0_expanded_f[0]}} & btb_bank0_rd_data_way0_f[BTB_DWIDTH - 1:0]) | ({17 + pt[2139-:9] {tag_match_way1_expanded_f[0]}} & btb_bank0_rd_data_way1_f[BTB_DWIDTH - 1:0]);
			assign btb_bank0e_rd_data_p1_f[BTB_DWIDTH - 1:0] = ({17 + pt[2139-:9] {tag_match_way0_expanded_p1_f[0]}} & btb_bank0_rd_data_way0_p1_f[BTB_DWIDTH - 1:0]) | ({17 + pt[2139-:9] {tag_match_way1_expanded_p1_f[0]}} & btb_bank0_rd_data_way1_p1_f[BTB_DWIDTH - 1:0]);
			wire [BTB_DWIDTH:1] sv2v_tmp_F09CF;
			assign sv2v_tmp_F09CF = ({17 + pt[2139-:9] {fetch_start_f[0]}} & btb_bank0e_rd_data_f[BTB_DWIDTH - 1:0]) | ({17 + pt[2139-:9] {fetch_start_f[1]}} & btb_bank0o_rd_data_f[BTB_DWIDTH - 1:0]);
			always @(*) btb_vbank0_rd_data_f[BTB_DWIDTH - 1:0] = sv2v_tmp_F09CF;
			wire [BTB_DWIDTH:1] sv2v_tmp_BEF15;
			assign sv2v_tmp_BEF15 = ({17 + pt[2139-:9] {fetch_start_f[0]}} & btb_bank0o_rd_data_f[BTB_DWIDTH - 1:0]) | ({17 + pt[2139-:9] {fetch_start_f[1]}} & btb_bank0e_rd_data_p1_f[BTB_DWIDTH - 1:0]);
			always @(*) btb_vbank1_rd_data_f[BTB_DWIDTH - 1:0] = sv2v_tmp_BEF15;
			assign way_raw[1:0] = tag_match_vway1_expanded_f[1:0] | (~vwayhit_f[1:0] & btb_vlru_rd_f[1:0]);
			assign mp_wrindex_dec[LRU_SIZE - 1:0] = {{LRU_SIZE - 1 {1'b0}}, 1'b1} << exu_mp_addr[pt[2172-:9]:pt[2163-:6]];
			assign fetch_wrindex_dec[LRU_SIZE - 1:0] = {{LRU_SIZE - 1 {1'b0}}, 1'b1} << btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]];
			assign fetch_wrindex_p1_dec[LRU_SIZE - 1:0] = {{LRU_SIZE - 1 {1'b0}}, 1'b1} << btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]];
			assign mp_wrlru_b0[LRU_SIZE - 1:0] = mp_wrindex_dec[LRU_SIZE - 1:0] & {LRU_SIZE {exu_mp_valid}};
			assign btb_lru_b0_hold[LRU_SIZE - 1:0] = ~mp_wrlru_b0[LRU_SIZE - 1:0] & ~fetch_wrlru_b0[LRU_SIZE - 1:0];
			assign use_mp_way = fetch_mp_collision_f;
			assign use_mp_way_p1 = fetch_mp_collision_p1_f;
			assign lru_update_valid_f = ((vwayhit_f[0] | vwayhit_f[1]) & ifc_fetch_req_f) & ~leak_one_f;
			assign fetch_wrlru_b0[LRU_SIZE - 1:0] = fetch_wrindex_dec[LRU_SIZE - 1:0] & {LRU_SIZE {lru_update_valid_f}};
			assign fetch_wrlru_p1_b0[LRU_SIZE - 1:0] = fetch_wrindex_p1_dec[LRU_SIZE - 1:0] & {LRU_SIZE {lru_update_valid_f}};
			assign btb_lru_b0_ns[LRU_SIZE - 1:0] = (((btb_lru_b0_hold[LRU_SIZE - 1:0] & btb_lru_b0_f[LRU_SIZE - 1:0]) | (mp_wrlru_b0[LRU_SIZE - 1:0] & {LRU_SIZE {~exu_mp_way}})) | (fetch_wrlru_b0[LRU_SIZE - 1:0] & {LRU_SIZE {tag_match_way0_f}})) | (fetch_wrlru_p1_b0[LRU_SIZE - 1:0] & {LRU_SIZE {tag_match_way0_p1_f}});
			assign btb_lru_rd_f = (use_mp_way ? exu_mp_way_f : |(fetch_wrindex_dec[LRU_SIZE - 1:0] & btb_lru_b0_f[LRU_SIZE - 1:0]));
			assign btb_lru_rd_p1_f = (use_mp_way_p1 ? exu_mp_way_f : |(fetch_wrindex_p1_dec[LRU_SIZE - 1:0] & btb_lru_b0_f[LRU_SIZE - 1:0]));
			assign btb_vlru_rd_f[1:0] = ({2 {fetch_start_f[0]}} & {btb_lru_rd_f, btb_lru_rd_f}) | ({2 {fetch_start_f[1]}} & {btb_lru_rd_p1_f, btb_lru_rd_f});
			assign tag_match_vway1_expanded_f[1:0] = ({2 {fetch_start_f[0]}} & {tag_match_way1_expanded_f[1:0]}) | ({2 {fetch_start_f[1]}} & {tag_match_way1_expanded_p1_f[0], tag_match_way1_expanded_f[1]});
			rvdffe #(.WIDTH(LRU_SIZE)) btb_lru_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(ifc_fetch_req_f | exu_mp_valid),
				.din(btb_lru_b0_ns[LRU_SIZE - 1:0]),
				.dout(btb_lru_b0_f[LRU_SIZE - 1:0])
			);
		end
	endgenerate
	wire eoc_near;
	wire eoc_mask;
	assign eoc_near = &ifc_fetch_addr_f[pt[1182-:8]:3];
	assign eoc_mask = ~eoc_near | |(~ifc_fetch_addr_f[2:1]);
	wire [16:1] btb_sel_data_f;
	assign btb_rd_tgt_f[11:0] = btb_sel_data_f[16:5];
	assign btb_rd_pc4_f = btb_sel_data_f[4];
	assign btb_rd_call_f = btb_sel_data_f[2];
	assign btb_rd_ret_f = btb_sel_data_f[1];
	assign btb_sel_data_f[16:1] = ({16 {btb_sel_f[1]}} & btb_vbank1_rd_data_f[16:1]) | ({16 {btb_sel_f[0]}} & btb_vbank0_rd_data_f[16:1]);
	wire [1:0] hist0_raw;
	wire [1:0] hist1_raw;
	wire [1:0] pc4_raw;
	wire [1:0] pret_raw;
	assign ifu_bp_hit_taken_f = ((|(vwayhit_f[1:0] & hist1_raw[1:0]) & ifc_fetch_req_f) & ~leak_one_f_d1) & ~dec_tlu_bpred_disable;
	assign bht_force_taken_f[1:0] = {btb_vbank1_rd_data_f[CALL] | btb_vbank1_rd_data_f[RET], btb_vbank0_rd_data_f[CALL] | btb_vbank0_rd_data_f[RET]};
	assign bht_valid_f[1:0] = vwayhit_f[1:0];
	assign bht_vbank0_rd_data_f[1:0] = ({2 {fetch_start_f[0]}} & bht_bank0_rd_data_f[1:0]) | ({2 {fetch_start_f[1]}} & bht_bank1_rd_data_f[1:0]);
	assign bht_vbank1_rd_data_f[1:0] = ({2 {fetch_start_f[0]}} & bht_bank1_rd_data_f[1:0]) | ({2 {fetch_start_f[1]}} & bht_bank0_rd_data_p1_f[1:0]);
	assign bht_dir_f[1:0] = {(bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]) & bht_valid_f[1], (bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]) & bht_valid_f[0]};
	assign ifu_bp_inst_mask_f = (ifu_bp_hit_taken_f & btb_sel_f[1]) | ~ifu_bp_hit_taken_f;
	assign hist1_raw[1:0] = bht_force_taken_f[1:0] | {bht_vbank1_rd_data_f[1], bht_vbank0_rd_data_f[1]};
	assign hist0_raw[1:0] = {bht_vbank1_rd_data_f[0], bht_vbank0_rd_data_f[0]};
	assign pc4_raw[1:0] = {vwayhit_f[1] & btb_vbank1_rd_data_f[PC4], vwayhit_f[0] & btb_vbank0_rd_data_f[PC4]};
	assign pret_raw[1:0] = {(vwayhit_f[1] & ~btb_vbank1_rd_data_f[CALL]) & btb_vbank1_rd_data_f[RET], (vwayhit_f[0] & ~btb_vbank0_rd_data_f[CALL]) & btb_vbank0_rd_data_f[RET]};
	function [1:0] countones;
		input [1:0] valid;
		countones[1:0] = {2'b00, valid[1]} + {2'b00, valid[0]};
	endfunction
	assign num_valids[1:0] = countones(bht_valid_f[1:0]);
	assign final_h = |(btb_sel_f[1:0] & bht_dir_f[1:0]);
	assign merged_ghr[pt[2236-:8] - 1:0] = (({pt[2236-:8] {num_valids[1:0] == 2'h2}} & {fghr[pt[2236-:8] - 3:0], 1'b0, final_h}) | ({pt[2236-:8] {num_valids[1:0] == 2'h1}} & {fghr[pt[2236-:8] - 2:0], final_h})) | ({pt[2236-:8] {num_valids[1:0] == 2'h0}} & {fghr[pt[2236-:8] - 1:0]});
	wire [pt[2236-:8] - 1:0] exu_flush_ghr;
	assign exu_flush_ghr[pt[2236-:8] - 1:0] = exu_mp_fghr[pt[2236-:8] - 1:0];
	assign fghr_ns[pt[2236-:8] - 1:0] = (({pt[2236-:8] {exu_flush_final_d1}} & exu_flush_ghr[pt[2236-:8] - 1:0]) | ({pt[2236-:8] {((~exu_flush_final_d1 & ifc_fetch_req_f) & ic_hit_f) & ~leak_one_f_d1}} & merged_ghr[pt[2236-:8] - 1:0])) | ({pt[2236-:8] {~exu_flush_final_d1 & ~((ifc_fetch_req_f & ic_hit_f) & ~leak_one_f_d1)}} & fghr[pt[2236-:8] - 1:0]);
	rvdffie #(
		.WIDTH(pt[2236-:8] + 3),
		.OVERRIDE(1)
	) fetchghr(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din({exu_flush_final, exu_mp_way, leak_one_f, fghr_ns[pt[2236-:8] - 1:0]}),
		.dout({exu_flush_final_d1, exu_mp_way_f, leak_one_f_d1, fghr[pt[2236-:8] - 1:0]})
	);
	assign ifu_bp_fghr_f[pt[2236-:8] - 1:0] = fghr[pt[2236-:8] - 1:0];
	assign ifu_bp_way_f[1:0] = way_raw[1:0];
	assign ifu_bp_hist1_f[1:0] = hist1_raw[1:0];
	assign ifu_bp_hist0_f[1:0] = hist0_raw[1:0];
	assign ifu_bp_pc4_f[1:0] = pc4_raw[1:0];
	assign ifu_bp_valid_f[1:0] = vwayhit_f[1:0] & ~{2 {dec_tlu_bpred_disable}};
	assign ifu_bp_ret_f[1:0] = pret_raw[1:0];
	wire [1:0] bloc_f;
	wire use_fa_plus;
	assign bloc_f[1] = (bht_dir_f[0] & ~fetch_start_f[0]) | (~bht_dir_f[0] & fetch_start_f[0]);
	assign bloc_f[0] = (bht_dir_f[0] & fetch_start_f[0]) | (~bht_dir_f[0] & ~fetch_start_f[0]);
	assign use_fa_plus = (~bht_dir_f[0] & ~fetch_start_f[0]) & ~btb_rd_pc4_f;
	assign btb_fg_crossing_f = (fetch_start_f[0] & btb_sel_f[0]) & btb_rd_pc4_f;
	assign bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f;
	wire [31:2] adder_pc_in_f;
	wire [31:2] ifc_fetch_adder_prior;
	rvdfflie #(
		.WIDTH(30),
		.LEFT(19)
	) faddrf_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((ifc_fetch_req_f & ~ifu_bp_hit_taken_f) & ic_hit_f),
		.din(ifc_fetch_addr_f[31:2]),
		.dout(ifc_fetch_adder_prior[31:2])
	);
	assign ifu_bp_poffset_f[11:0] = btb_rd_tgt_f[11:0];
	assign adder_pc_in_f[31:2] = (({30 {use_fa_plus}} & fetch_addr_p1_f[31:2]) | ({30 {btb_fg_crossing_f}} & ifc_fetch_adder_prior[31:2])) | ({30 {~btb_fg_crossing_f & ~use_fa_plus}} & ifc_fetch_addr_f[31:2]);
	rvbradder predtgt_addr(
		.pc({adder_pc_in_f[31:2], bp_total_branch_offset_f}),
		.offset(btb_rd_tgt_f[11:0]),
		.dout(bp_btb_target_adder_f[31:1])
	);
	assign ifu_bp_btb_target_f[31:1] = ({31 {((btb_rd_ret_f & ~btb_rd_call_f) & rets_out[0]) & ifu_bp_hit_taken_f}} & rets_out[31-:31]) | ({31 {~((btb_rd_ret_f & ~btb_rd_call_f) & rets_out[0]) & ifu_bp_hit_taken_f}} & bp_btb_target_adder_f[31:1]);
	rvbradder rs_addr(
		.pc({adder_pc_in_f[31:2], bp_total_branch_offset_f}),
		.offset({11'b00000000000, ~btb_rd_pc4_f}),
		.dout(bp_rs_call_target_f[31:1])
	);
	assign rs_push = (btb_rd_call_f & ~btb_rd_ret_f) & ifu_bp_hit_taken_f;
	assign rs_pop = (btb_rd_ret_f & ~btb_rd_call_f) & ifu_bp_hit_taken_f;
	assign rs_hold = ~rs_push & ~rs_pop;
	assign rets_in[31-:32] = ({32 {rs_push}} & {bp_rs_call_target_f[31:1], 1'b1}) | ({32 {rs_pop}} & rets_out[63-:32]);
	assign rsenable[0] = ~rs_hold;
	generate
		for (i = 0; i < pt[31-:8]; i = i + 1) begin : retstack
			if (i == (pt[31-:8] - 1)) begin
				assign rets_in[(i * 32) + 31-:32] = rets_out[((i - 1) * 32) + 31-:32];
				assign rsenable[i] = rs_push;
			end
			else if (i > 0) begin
				assign rets_in[(i * 32) + 31-:32] = ({32 {rs_push}} & rets_out[((i - 1) * 32) + 31-:32]) | ({32 {rs_pop}} & rets_out[((i + 1) * 32) + 31-:32]);
				assign rsenable[i] = rs_push | rs_pop;
			end
			rvdffe #(.WIDTH(32)) rets_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(rsenable[i]),
				.din(rets_in[(i * 32) + 31-:32]),
				.dout(rets_out[(i * 32) + 31-:32])
			);
		end
	endgenerate
	assign dec_tlu_error_wb = dec_tlu_br0_start_error_wb | dec_tlu_br0_error_wb;
	assign btb_error_addr_wb[pt[2172-:9]:pt[2163-:6]] = dec_tlu_br0_addr_wb[pt[2172-:9]:pt[2163-:6]];
	assign dec_tlu_way_wb = dec_tlu_br0_way_wb;
	assign btb_valid = exu_mp_valid & ~dec_tlu_error_wb;
	assign btb_wr_tag[pt[2139-:9] - 1:0] = exu_mp_btag[pt[2139-:9] - 1:0];
	generate
		if (!pt[2120-:5]) begin
			if (pt[2144-:5]) begin : btbfold
				eb1_btb_tag_hash_fold #(.pt(pt)) rdtagf(
					.hash(fetch_rd_tag_f[pt[2139-:9] - 1:0]),
					.pc({ifc_fetch_addr_f[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]})
				);
				eb1_btb_tag_hash_fold #(.pt(pt)) rdtagp1f(
					.hash(fetch_rd_tag_p1_f[pt[2139-:9] - 1:0]),
					.pc({fetch_addr_p1_f[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]})
				);
			end
			else begin
				eb1_btb_tag_hash #(.pt(pt)) rdtagf(
					.hash(fetch_rd_tag_f[pt[2139-:9] - 1:0]),
					.pc({ifc_fetch_addr_f[((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]})
				);
				eb1_btb_tag_hash #(.pt(pt)) rdtagp1f(
					.hash(fetch_rd_tag_p1_f[pt[2139-:9] - 1:0]),
					.pc({fetch_addr_p1_f[((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1]})
				);
			end
			assign btb_wr_en_way0 = {(~exu_mp_way & exu_mp_valid_write) & ~dec_tlu_error_wb} | {~dec_tlu_way_wb & dec_tlu_error_wb};
			assign btb_wr_en_way1 = {(exu_mp_way & exu_mp_valid_write) & ~dec_tlu_error_wb} | {dec_tlu_way_wb & dec_tlu_error_wb};
			assign btb_wr_addr[pt[2172-:9]:pt[2163-:6]] = (dec_tlu_error_wb ? btb_error_addr_wb[pt[2172-:9]:pt[2163-:6]] : exu_mp_addr[pt[2172-:9]:pt[2163-:6]]);
			assign vwayhit_f[1:0] = (({2 {fetch_start_f[0]}} & {wayhit_f[1:0]}) | ({2 {fetch_start_f[1]}} & {wayhit_p1_f[0], wayhit_f[1]})) & {eoc_mask, 1'b1};
		end
	endgenerate
	assign btb_wr_data[BTB_DWIDTH - 1:0] = {btb_wr_tag[pt[2139-:9] - 1:0], exu_mp_tgt[pt[2047-:9] - 1:0], exu_mp_pc4, exu_mp_boffset, exu_mp_call | exu_mp_ja, exu_mp_ret | exu_mp_ja, btb_valid};
	assign exu_mp_valid_write = (exu_mp_valid & exu_mp_ataken) & ~exu_mp_pkt[37];
	wire [1:0] bht_wr_data0;
	wire [1:0] bht_wr_data2;
	wire [1:0] bht_wr_en0;
	wire [1:0] bht_wr_en2;
	assign middle_of_bank = exu_mp_pc4 ^ exu_mp_boffset;
	assign bht_wr_en0[1:0] = {2 {((exu_mp_valid & ~exu_mp_call) & ~exu_mp_ret) & ~exu_mp_ja}} & {middle_of_bank, ~middle_of_bank};
	assign bht_wr_en2[1:0] = {2 {dec_tlu_br0_v_wb}} & {dec_tlu_br0_middle_wb, ~dec_tlu_br0_middle_wb};
	assign bht_wr_data0[1:0] = exu_mp_hist[1:0];
	assign bht_wr_data2[1:0] = dec_tlu_br0_hist_wb[1:0];
	wire [pt[2270-:8]:pt[2262-:6]] bht_rd_addr_f;
	wire [pt[2270-:8]:pt[2262-:6]] bht_rd_addr_p1_f;
	wire [pt[2270-:8]:pt[2262-:6]] bht_wr_addr0;
	wire [pt[2270-:8]:pt[2262-:6]] bht_wr_addr2;
	wire [pt[2270-:8]:pt[2262-:6]] mp_hashed;
	wire [pt[2270-:8]:pt[2262-:6]] br0_hashed_wb;
	wire [pt[2270-:8]:pt[2262-:6]] bht_rd_addr_hashed_f;
	wire [pt[2270-:8]:pt[2262-:6]] bht_rd_addr_hashed_p1_f;
	eb1_btb_ghr_hash #(.pt(pt)) mpghrhs(
		.hashin(exu_mp_addr[pt[2172-:9]:pt[2163-:6]]),
		.ghr(exu_mp_eghr[pt[2236-:8] - 1:0]),
		.hash(mp_hashed[pt[2270-:8]:pt[2262-:6]])
	);
	eb1_btb_ghr_hash #(.pt(pt)) br0ghrhs(
		.hashin(dec_tlu_br0_addr_wb[pt[2172-:9]:pt[2163-:6]]),
		.ghr(exu_i0_br_fghr_wb[pt[2236-:8] - 1:0]),
		.hash(br0_hashed_wb[pt[2270-:8]:pt[2262-:6]])
	);
	eb1_btb_ghr_hash #(.pt(pt)) fghrhs(
		.hashin(btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]]),
		.ghr(fghr[pt[2236-:8] - 1:0]),
		.hash(bht_rd_addr_hashed_f[pt[2270-:8]:pt[2262-:6]])
	);
	eb1_btb_ghr_hash #(.pt(pt)) fghrhs_p1(
		.hashin(btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]]),
		.ghr(fghr[pt[2236-:8] - 1:0]),
		.hash(bht_rd_addr_hashed_p1_f[pt[2270-:8]:pt[2262-:6]])
	);
	assign bht_wr_addr0[pt[2270-:8]:pt[2262-:6]] = mp_hashed[pt[2270-:8]:pt[2262-:6]];
	assign bht_wr_addr2[pt[2270-:8]:pt[2262-:6]] = br0_hashed_wb[pt[2270-:8]:pt[2262-:6]];
	assign bht_rd_addr_f[pt[2270-:8]:pt[2262-:6]] = bht_rd_addr_hashed_f[pt[2270-:8]:pt[2262-:6]];
	assign bht_rd_addr_p1_f[pt[2270-:8]:pt[2262-:6]] = bht_rd_addr_hashed_p1_f[pt[2270-:8]:pt[2262-:6]];
	generate
		if (!pt[2120-:5]) begin
			for (j = 0; j < LRU_SIZE; j = j + 1) begin : BTB_FLOPS
				rvdffe #(.WIDTH(17 + pt[2139-:9])) btb_bank0_way0(
					.clk(clk),
					.rst_l(rst_l),
					.scan_mode(scan_mode),
					.en((btb_wr_addr[pt[2172-:9]:pt[2163-:6]] == j) & btb_wr_en_way0),
					.din(btb_wr_data[BTB_DWIDTH - 1:0]),
					.dout(btb_bank0_rd_data_way0_out[j * BTB_DWIDTH+:BTB_DWIDTH])
				);
				rvdffe #(.WIDTH(17 + pt[2139-:9])) btb_bank0_way1(
					.clk(clk),
					.rst_l(rst_l),
					.scan_mode(scan_mode),
					.en((btb_wr_addr[pt[2172-:9]:pt[2163-:6]] == j) & btb_wr_en_way1),
					.din(btb_wr_data[BTB_DWIDTH - 1:0]),
					.dout(btb_bank0_rd_data_way1_out[j * BTB_DWIDTH+:BTB_DWIDTH])
				);
			end
			function automatic signed [((pt[2172-:9] - pt[2163-:6]) >= 0 ? (pt[2172-:9] - pt[2163-:6]) + 1 : 1 - (pt[2172-:9] - pt[2163-:6])) - 1:0] sv2v_cast_C4842_signed;
				input reg signed [((pt[2172-:9] - pt[2163-:6]) >= 0 ? (pt[2172-:9] - pt[2163-:6]) + 1 : 1 - (pt[2172-:9] - pt[2163-:6])) - 1:0] inp;
				sv2v_cast_C4842_signed = inp;
			endfunction
			always @(*) begin : BTB_rd_mux
				btb_bank0_rd_data_way0_f[BTB_DWIDTH - 1:0] = {BTB_DWIDTH {1'sb0}};
				btb_bank0_rd_data_way1_f[BTB_DWIDTH - 1:0] = {BTB_DWIDTH {1'sb0}};
				btb_bank0_rd_data_way0_p1_f[BTB_DWIDTH - 1:0] = {BTB_DWIDTH {1'sb0}};
				btb_bank0_rd_data_way1_p1_f[BTB_DWIDTH - 1:0] = {BTB_DWIDTH {1'sb0}};
				begin : sv2v_autoblock_43
					reg signed [31:0] j;
					for (j = 0; j < LRU_SIZE; j = j + 1)
						if (btb_rd_addr_f[pt[2172-:9]:pt[2163-:6]] == sv2v_cast_C4842_signed(j)) begin
							btb_bank0_rd_data_way0_f[BTB_DWIDTH - 1:0] = btb_bank0_rd_data_way0_out[j * BTB_DWIDTH+:BTB_DWIDTH];
							btb_bank0_rd_data_way1_f[BTB_DWIDTH - 1:0] = btb_bank0_rd_data_way1_out[j * BTB_DWIDTH+:BTB_DWIDTH];
						end
				end
				begin : sv2v_autoblock_44
					reg signed [31:0] j;
					for (j = 0; j < LRU_SIZE; j = j + 1)
						if (btb_rd_addr_p1_f[pt[2172-:9]:pt[2163-:6]] == sv2v_cast_C4842_signed(j)) begin
							btb_bank0_rd_data_way0_p1_f[BTB_DWIDTH - 1:0] = btb_bank0_rd_data_way0_out[j * BTB_DWIDTH+:BTB_DWIDTH];
							btb_bank0_rd_data_way1_p1_f[BTB_DWIDTH - 1:0] = btb_bank0_rd_data_way1_out[j * BTB_DWIDTH+:BTB_DWIDTH];
						end
				end
			end
		end
	endgenerate
	generate
		if (pt[2120-:5]) begin : fa
			reg found1;
			reg hit0;
			reg hit1;
			wire btb_used_reset;
			wire write_used;
			reg [$clog2(pt[2061-:14]) - 1:0] btb_fa_wr_addr0;
			reg [$clog2(pt[2061-:14]) - 1:0] hit0_index;
			reg [$clog2(pt[2061-:14]) - 1:0] hit1_index;
			reg [pt[2061-:14] - 1:0] btb_tag_hit;
			reg [pt[2061-:14] - 1:0] btb_offset_0;
			reg [pt[2061-:14] - 1:0] btb_offset_1;
			wire [pt[2061-:14] - 1:0] btb_used_ns;
			wire [pt[2061-:14] - 1:0] btb_used;
			wire [pt[2061-:14] - 1:0] wr0_en;
			reg [pt[2061-:14] - 1:0] btb_upper_hit;
			wire [(pt[2061-:14] * BTB_DWIDTH) - 1:0] btbdata;
			wire [FA_CMP_LOWER - 1:1] ifc_fetch_addr_p1_f;
			assign ifc_fetch_addr_p1_f[FA_CMP_LOWER - 1:1] = ifc_fetch_addr_f[FA_CMP_LOWER - 1:1] + 1'b1;
			assign fetch_mp_collision_f = (((exu_mp_btag[pt[2139-:9] - 1:0] == ifc_fetch_addr_f[31:1]) & exu_mp_valid) & ifc_fetch_req_f) & ~exu_mp_pkt[32];
			assign fetch_mp_collision_p1_f = (((exu_mp_btag[pt[2139-:9] - 1:0] == {ifc_fetch_addr_f[31:FA_CMP_LOWER], ifc_fetch_addr_p1_f[FA_CMP_LOWER - 1:1]}) & exu_mp_valid) & ifc_fetch_req_f) & ~exu_mp_pkt[32];
			function automatic signed [(BTB_FA_INDEX >= 0 ? BTB_FA_INDEX + 1 : 1 - BTB_FA_INDEX) - 1:0] sv2v_cast_50CAB_signed;
				input reg signed [(BTB_FA_INDEX >= 0 ? BTB_FA_INDEX + 1 : 1 - BTB_FA_INDEX) - 1:0] inp;
				sv2v_cast_50CAB_signed = inp;
			endfunction
			always @(*) begin
				btb_vbank0_rd_data_f = {BTB_DWIDTH {1'sb0}};
				btb_vbank1_rd_data_f = {BTB_DWIDTH {1'sb0}};
				btb_tag_hit = {pt[2061-:14] {1'sb0}};
				btb_upper_hit = {pt[2061-:14] {1'sb0}};
				btb_offset_0 = {pt[2061-:14] {1'sb0}};
				btb_offset_1 = {pt[2061-:14] {1'sb0}};
				found1 = 1'b0;
				hit0 = 1'b0;
				hit1 = 1'b0;
				hit0_index = {$clog2(pt[2061-:14]) {1'sb0}};
				hit1_index = {$clog2(pt[2061-:14]) {1'sb0}};
				btb_fa_wr_addr0 = {$clog2(pt[2061-:14]) {1'sb0}};
				begin : sv2v_autoblock_45
					reg signed [31:0] i;
					for (i = 0; i < pt[2061-:14]; i = i + 1)
						begin
							btb_upper_hit[i] = ((btbdata[(i * BTB_DWIDTH) + (BTB_DWIDTH_TOP >= FA_TAG_END_UPPER ? BTB_DWIDTH_TOP : (BTB_DWIDTH_TOP + (BTB_DWIDTH_TOP >= FA_TAG_END_UPPER ? (BTB_DWIDTH_TOP - FA_TAG_END_UPPER) + 1 : (FA_TAG_END_UPPER - BTB_DWIDTH_TOP) + 1)) - 1)-:(BTB_DWIDTH_TOP >= FA_TAG_END_UPPER ? (BTB_DWIDTH_TOP - FA_TAG_END_UPPER) + 1 : (FA_TAG_END_UPPER - BTB_DWIDTH_TOP) + 1)] == ifc_fetch_addr_f[31:FA_CMP_LOWER]) & btbdata[i * BTB_DWIDTH]) & ~wr0_en[i];
							btb_offset_0[i] = (btbdata[(i * BTB_DWIDTH) + (FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? FA_TAG_START_LOWER : (FA_TAG_START_LOWER + (FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? (FA_TAG_START_LOWER - FA_TAG_END_LOWER) + 1 : (FA_TAG_END_LOWER - FA_TAG_START_LOWER) + 1)) - 1)-:(FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? (FA_TAG_START_LOWER - FA_TAG_END_LOWER) + 1 : (FA_TAG_END_LOWER - FA_TAG_START_LOWER) + 1)] == ifc_fetch_addr_f[FA_CMP_LOWER - 1:1]) & btb_upper_hit[i];
							btb_offset_1[i] = (btbdata[(i * BTB_DWIDTH) + (FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? FA_TAG_START_LOWER : (FA_TAG_START_LOWER + (FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? (FA_TAG_START_LOWER - FA_TAG_END_LOWER) + 1 : (FA_TAG_END_LOWER - FA_TAG_START_LOWER) + 1)) - 1)-:(FA_TAG_START_LOWER >= FA_TAG_END_LOWER ? (FA_TAG_START_LOWER - FA_TAG_END_LOWER) + 1 : (FA_TAG_END_LOWER - FA_TAG_START_LOWER) + 1)] == ifc_fetch_addr_p1_f[FA_CMP_LOWER - 1:1]) & btb_upper_hit[i];
							if (~hit0)
								if (btb_offset_0[i]) begin
									hit0_index[BTB_FA_INDEX:0] = sv2v_cast_50CAB_signed(i);
									hit0 = 1'b1;
								end
							if (~hit1)
								if (btb_offset_1[i]) begin
									hit1_index[BTB_FA_INDEX:0] = sv2v_cast_50CAB_signed(i);
									hit1 = 1'b1;
								end
							if (btb_offset_0[i] == 1'b1)
								btb_vbank0_rd_data_f[BTB_DWIDTH - 1:0] = (fetch_mp_collision_f ? btb_wr_data : btbdata[i * BTB_DWIDTH+:BTB_DWIDTH]);
							if (btb_offset_1[i] == 1'b1)
								btb_vbank1_rd_data_f[BTB_DWIDTH - 1:0] = (fetch_mp_collision_p1_f ? btb_wr_data : btbdata[i * BTB_DWIDTH+:BTB_DWIDTH]);
							if (~found1)
								if (~btb_used[i]) begin
									btb_fa_wr_addr0[BTB_FA_INDEX:0] = i[BTB_FA_INDEX:0];
									found1 = 1'b1;
								end
						end
				end
			end
			assign vwayhit_f[1:0] = {hit1, hit0} & {eoc_mask, 1'b1};
			assign way_raw[1:0] = vwayhit_f[1:0] | {fetch_mp_collision_p1_f, fetch_mp_collision_f};
			for (j = 0; j < pt[2061-:14]; j = j + 1) begin : BTB_FAFLOPS
				assign wr0_en[j] = ((btb_fa_wr_addr0[BTB_FA_INDEX:0] == j) & (exu_mp_valid_write & ~exu_mp_pkt[32])) | ((dec_fa_error_index == j) & dec_tlu_error_wb);
				rvdffe #(.WIDTH(BTB_DWIDTH)) btb_fa(
					.rst_l(rst_l),
					.scan_mode(scan_mode),
					.clk(clk),
					.en(wr0_en[j]),
					.din(btb_wr_data[BTB_DWIDTH - 1:0]),
					.dout(btbdata[j * BTB_DWIDTH+:BTB_DWIDTH])
				);
			end
			assign ifu_bp_fa_index_f[$clog2(pt[2061-:14])+:$clog2(pt[2061-:14])] = (hit1 ? hit1_index : {$clog2(pt[2061-:14]) {1'sb0}});
			assign ifu_bp_fa_index_f[0+:$clog2(pt[2061-:14])] = (hit0 ? hit0_index : {$clog2(pt[2061-:14]) {1'sb0}});
			assign btb_used_reset = &btb_used[pt[2061-:14] - 1:0];
			assign btb_used_ns[pt[2061-:14] - 1:0] = ((((({pt[2061-:14] {vwayhit_f[1]}} & (32'b00000000000000000000000000000001 << hit1_index[BTB_FA_INDEX:0])) | ({pt[2061-:14] {vwayhit_f[0]}} & (32'b00000000000000000000000000000001 << hit0_index[BTB_FA_INDEX:0]))) | ({pt[2061-:14] {(exu_mp_valid_write & ~exu_mp_pkt[32]) & ~dec_tlu_error_wb}} & (32'b00000000000000000000000000000001 << btb_fa_wr_addr0[BTB_FA_INDEX:0]))) | ({pt[2061-:14] {btb_used_reset}} & {pt[2061-:14] {1'b0}})) | ({pt[2061-:14] {~btb_used_reset & dec_tlu_error_wb}} & (btb_used[pt[2061-:14] - 1:0] & ~(32'b00000000000000000000000000000001 << dec_fa_error_index[BTB_FA_INDEX:0])))) | (~{pt[2061-:14] {btb_used_reset | dec_tlu_error_wb}} & btb_used[pt[2061-:14] - 1:0]);
			assign write_used = ((btb_used_reset | ifu_bp_hit_taken_f) | exu_mp_valid_write) | dec_tlu_error_wb;
			rvdffe #(.WIDTH(pt[2061-:14])) btb_usedf(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(write_used),
				.din(btb_used_ns[pt[2061-:14] - 1:0]),
				.dout(btb_used[pt[2061-:14] - 1:0])
			);
		end
	endgenerate
	wire [(((2 * (pt[2256-:15] / NUM_BHT_LOOP)) * NUM_BHT_LOOP) * 2) - 1:0] bht_bank_wr_data;
	wire [((2 * pt[2256-:15]) * 2) - 1:0] bht_bank_rd_data_out;
	wire [(2 * (pt[2256-:15] / NUM_BHT_LOOP)) - 1:0] bht_bank_clken;
	wire [(2 * (pt[2256-:15] / NUM_BHT_LOOP)) - 1:0] bht_bank_clk;
	wire [((2 * (pt[2256-:15] / NUM_BHT_LOOP)) * NUM_BHT_LOOP) - 1:0] bht_bank_sel;
	generate
		for (i = 0; i < 2; i = i + 1) begin : BANKS
			genvar k;
			for (k = 0; k < (pt[2256-:15] / NUM_BHT_LOOP); k = k + 1) begin : BHT_CLK_GROUP
				assign bht_bank_clken[(i * (pt[2256-:15] / NUM_BHT_LOOP)) + k] = (bht_wr_en0[i] & ((bht_wr_addr0[pt[2270-:8]:NUM_BHT_LOOP_OUTER_LO] == k) | BHT_NO_ADDR_MATCH)) | (bht_wr_en2[i] & ((bht_wr_addr2[pt[2270-:8]:NUM_BHT_LOOP_OUTER_LO] == k) | BHT_NO_ADDR_MATCH));
				rvclkhdr bht_bank_grp_cgc(
					.en(bht_bank_clken[(i * (pt[2256-:15] / NUM_BHT_LOOP)) + k]),
					.l1clk(bht_bank_clk[(i * (pt[2256-:15] / NUM_BHT_LOOP)) + k]),
					.clk(clk),
					.scan_mode(scan_mode)
				);
				for (j = 0; j < NUM_BHT_LOOP; j = j + 1) begin : BHT_FLOPS
					assign bht_bank_sel[(((i * (pt[2256-:15] / NUM_BHT_LOOP)) + k) * NUM_BHT_LOOP) + j] = ((bht_wr_en0[i] & (bht_wr_addr0[NUM_BHT_LOOP_INNER_HI:pt[2262-:6]] == j)) & ((bht_wr_addr0[pt[2270-:8]:NUM_BHT_LOOP_OUTER_LO] == k) | BHT_NO_ADDR_MATCH)) | ((bht_wr_en2[i] & (bht_wr_addr2[NUM_BHT_LOOP_INNER_HI:pt[2262-:6]] == j)) & ((bht_wr_addr2[pt[2270-:8]:NUM_BHT_LOOP_OUTER_LO] == k) | BHT_NO_ADDR_MATCH));
					assign bht_bank_wr_data[((((i * (pt[2256-:15] / NUM_BHT_LOOP)) + k) * NUM_BHT_LOOP) + j) * 2+:2] = ((bht_wr_en2[i] & (bht_wr_addr2[NUM_BHT_LOOP_INNER_HI:pt[2262-:6]] == j)) & ((bht_wr_addr2[pt[2270-:8]:NUM_BHT_LOOP_OUTER_LO] == k) | BHT_NO_ADDR_MATCH) ? bht_wr_data2[1:0] : bht_wr_data0[1:0]);
					rvdffs_fpga #(.WIDTH(2)) bht_bank(
						.rst_l(rst_l),
						.clk(bht_bank_clk[(i * (pt[2256-:15] / NUM_BHT_LOOP)) + k]),
						.en(bht_bank_sel[(((i * (pt[2256-:15] / NUM_BHT_LOOP)) + k) * NUM_BHT_LOOP) + j]),
						.rawclk(clk),
						.clken(bht_bank_sel[(((i * (pt[2256-:15] / NUM_BHT_LOOP)) + k) * NUM_BHT_LOOP) + j]),
						.din(bht_bank_wr_data[((((i * (pt[2256-:15] / NUM_BHT_LOOP)) + k) * NUM_BHT_LOOP) + j) * 2+:2]),
						.dout(bht_bank_rd_data_out[((i * pt[2256-:15]) + ((16 * k) + j)) * 2+:2])
					);
				end
			end
		end
	endgenerate
	function automatic signed [((pt[2270-:8] - pt[2262-:6]) >= 0 ? (pt[2270-:8] - pt[2262-:6]) + 1 : 1 - (pt[2270-:8] - pt[2262-:6])) - 1:0] sv2v_cast_AB44B_signed;
		input reg signed [((pt[2270-:8] - pt[2262-:6]) >= 0 ? (pt[2270-:8] - pt[2262-:6]) + 1 : 1 - (pt[2270-:8] - pt[2262-:6])) - 1:0] inp;
		sv2v_cast_AB44B_signed = inp;
	endfunction
	always @(*) begin : BHT_rd_mux
		bht_bank0_rd_data_f[1:0] = {2 {1'sb0}};
		bht_bank1_rd_data_f[1:0] = {2 {1'sb0}};
		bht_bank0_rd_data_p1_f[1:0] = {2 {1'sb0}};
		begin : sv2v_autoblock_46
			reg signed [31:0] j;
			for (j = 0; j < pt[2256-:15]; j = j + 1)
				begin
					if (bht_rd_addr_f[pt[2270-:8]:pt[2262-:6]] == sv2v_cast_AB44B_signed(j)) begin
						bht_bank0_rd_data_f[1:0] = bht_bank_rd_data_out[j * 2+:2];
						bht_bank1_rd_data_f[1:0] = bht_bank_rd_data_out[(pt[2256-:15] + j) * 2+:2];
					end
					if (bht_rd_addr_p1_f[pt[2270-:8]:pt[2262-:6]] == sv2v_cast_AB44B_signed(j))
						bht_bank0_rd_data_p1_f[1:0] = bht_bank_rd_data_out[j * 2+:2];
				end
		end
	end
endmodule
module eb1_ifu_compress_ctl (
	din,
	dout
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [15:0] din;
	output wire [31:0] dout;
	wire legal;
	wire [15:0] i;
	wire [31:0] o;
	wire [31:0] l1;
	wire [31:0] l2;
	wire [31:0] l3;
	assign i[15:0] = din[15:0];
	wire [4:0] rs2d;
	wire [4:0] rdd;
	wire [4:0] rdpd;
	wire [4:0] rs2pd;
	wire rdrd;
	wire rdrs1;
	wire rs2rs2;
	wire rdprd;
	wire rdprs1;
	wire rs2prs2;
	wire rs2prd;
	wire uimm9_2;
	wire ulwimm6_2;
	wire ulwspimm7_2;
	wire rdeq2;
	wire rdeq1;
	wire rs1eq2;
	wire sbroffset8_1;
	wire simm9_4;
	wire simm5_0;
	wire sjaloffset11_1;
	wire sluimm17_12;
	wire uimm5_0;
	wire uswimm6_2;
	wire uswspimm7_2;
	assign rs2d[4:0] = i[6:2];
	assign rdd[4:0] = i[11:7];
	assign rdpd[4:0] = {2'b01, i[9:7]};
	assign rs2pd[4:0] = {2'b01, i[4:2]};
	assign l1[6:0] = o[6:0];
	assign l1[11:7] = ((((o[11:7] | ({5 {rdrd}} & rdd[4:0])) | ({5 {rdprd}} & rdpd[4:0])) | ({5 {rs2prd}} & rs2pd[4:0])) | ({5 {rdeq1}} & 5'd1)) | ({5 {rdeq2}} & 5'd2);
	assign l1[14:12] = o[14:12];
	assign l1[19:15] = ((o[19:15] | ({5 {rdrs1}} & rdd[4:0])) | ({5 {rdprs1}} & rdpd[4:0])) | ({5 {rs1eq2}} & 5'd2);
	assign l1[24:20] = (o[24:20] | ({5 {rs2rs2}} & rs2d[4:0])) | ({5 {rs2prs2}} & rs2pd[4:0]);
	assign l1[31:25] = o[31:25];
	wire [5:0] simm5d;
	wire [9:2] uimm9d;
	wire [9:4] simm9d;
	wire [6:2] ulwimm6d;
	wire [7:2] ulwspimm7d;
	wire [5:0] uimm5d;
	wire [20:1] sjald;
	wire [31:12] sluimmd;
	assign simm5d[5:0] = {i[12], i[6:2]};
	assign uimm9d[9:2] = {i[10:7], i[12:11], i[5], i[6]};
	assign simm9d[9:4] = {i[12], i[4:3], i[5], i[2], i[6]};
	assign ulwimm6d[6:2] = {i[5], i[12:10], i[6]};
	assign ulwspimm7d[7:2] = {i[3:2], i[12], i[6:4]};
	assign uimm5d[5:0] = {i[12], i[6:2]};
	assign sjald[11:1] = {i[12], i[8], i[10:9], i[6], i[7], i[2], i[11], i[5:4], i[3]};
	assign sjald[20:12] = {9 {i[12]}};
	assign sluimmd[31:12] = {{15 {i[12]}}, i[6:2]};
	assign l2[31:20] = (((((((l1[31:20] | ({12 {simm5_0}} & {{7 {simm5d[5]}}, simm5d[4:0]})) | ({12 {uimm9_2}} & {2'b00, uimm9d[9:2], 2'b00})) | ({12 {simm9_4}} & {{3 {simm9d[9]}}, simm9d[8:4], 4'b0000})) | ({12 {ulwimm6_2}} & {5'b00000, ulwimm6d[6:2], 2'b00})) | ({12 {ulwspimm7_2}} & {4'b0000, ulwspimm7d[7:2], 2'b00})) | ({12 {uimm5_0}} & {6'b000000, uimm5d[5:0]})) | ({12 {sjaloffset11_1}} & {sjald[20], sjald[10:1], sjald[11]})) | ({12 {sluimm17_12}} & sluimmd[31:20]);
	assign l2[19:12] = (l1[19:12] | ({8 {sjaloffset11_1}} & sjald[19:12])) | ({8 {sluimm17_12}} & sluimmd[19:12]);
	assign l2[11:0] = l1[11:0];
	wire [8:1] sbr8d;
	wire [6:2] uswimm6d;
	wire [7:2] uswspimm7d;
	assign sbr8d[8:1] = {i[12], i[6], i[5], i[2], i[11], i[10], i[4], i[3]};
	assign uswimm6d[6:2] = {i[5], i[12:10], i[6]};
	assign uswspimm7d[7:2] = {i[8:7], i[12:9]};
	assign l3[31:25] = ((l2[31:25] | ({7 {sbroffset8_1}} & {{4 {sbr8d[8]}}, sbr8d[7:5]})) | ({7 {uswimm6_2}} & {5'b00000, uswimm6d[6:5]})) | ({7 {uswspimm7_2}} & {4'b0000, uswspimm7d[7:5]});
	assign l3[24:12] = l2[24:12];
	assign l3[11:7] = ((l2[11:7] | ({5 {sbroffset8_1}} & {sbr8d[4:1], sbr8d[8]})) | ({5 {uswimm6_2}} & {uswimm6d[4:2], 2'b00})) | ({5 {uswspimm7_2}} & {uswspimm7d[4:2], 2'b00});
	assign l3[6:0] = l2[6:0];
	assign dout[31:0] = l3[31:0] & {32 {legal}};
	assign rdrd = ((((((((((((!i[14] & i[6]) & i[1]) | (((!i[15] & i[14]) & i[11]) & i[0])) | ((!i[14] & i[5]) & i[1])) | (((!i[15] & i[14]) & i[10]) & i[0])) | ((!i[14] & i[4]) & i[1])) | (((!i[15] & i[14]) & i[9]) & i[0])) | ((!i[14] & i[3]) & i[1])) | (((!i[15] & i[14]) & !i[8]) & i[0])) | ((!i[14] & i[2]) & i[1])) | (((!i[15] & i[14]) & i[7]) & i[0])) | (!i[15] & i[1])) | ((!i[15] & !i[13]) & i[0]);
	assign rdrs1 = ((((((((((((((!i[14] & i[12]) & i[11]) & i[1]) | (((!i[14] & i[12]) & i[10]) & i[1])) | (((!i[14] & i[12]) & i[9]) & i[1])) | (((!i[14] & i[12]) & i[8]) & i[1])) | (((!i[14] & i[12]) & i[7]) & i[1])) | (((((((!i[14] & !i[12]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | (((!i[14] & i[12]) & i[6]) & i[1])) | (((!i[14] & i[12]) & i[5]) & i[1])) | (((!i[14] & i[12]) & i[4]) & i[1])) | (((!i[14] & i[12]) & i[3]) & i[1])) | (((!i[14] & i[12]) & i[2]) & i[1])) | (((!i[15] & !i[14]) & !i[13]) & i[0])) | ((!i[15] & !i[14]) & i[1]);
	assign rs2rs2 = ((((((i[15] & i[6]) & i[1]) | ((i[15] & i[5]) & i[1])) | ((i[15] & i[4]) & i[1])) | ((i[15] & i[3]) & i[1])) | ((i[15] & i[2]) & i[1])) | ((i[15] & i[14]) & i[1]);
	assign rdprd = ((i[15] & !i[14]) & !i[13]) & i[0];
	assign rdprs1 = (((i[15] & !i[13]) & i[0]) | ((i[15] & i[14]) & i[0])) | ((i[14] & !i[1]) & !i[0]);
	assign rs2prs2 = (((((i[15] & !i[14]) & !i[13]) & i[11]) & i[10]) & i[0]) | ((i[15] & !i[1]) & !i[0]);
	assign rs2prd = (!i[15] & !i[1]) & !i[0];
	assign uimm9_2 = (!i[14] & !i[1]) & !i[0];
	assign ulwimm6_2 = ((!i[15] & i[14]) & !i[1]) & !i[0];
	assign ulwspimm7_2 = (!i[15] & i[14]) & i[1];
	assign rdeq2 = ((((((!i[15] & i[14]) & i[13]) & !i[11]) & !i[10]) & !i[9]) & i[8]) & !i[7];
	assign rdeq1 = ((((((((((((!i[14] & i[12]) & i[11]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1]) | ((((((((!i[14] & i[12]) & i[10]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[9]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[8]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[7]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((!i[15] & !i[14]) & i[13]);
	assign rs1eq2 = ((((((((!i[15] & i[14]) & i[13]) & !i[11]) & !i[10]) & !i[9]) & i[8]) & !i[7]) | (i[14] & i[1])) | ((!i[14] & !i[1]) & !i[0]);
	assign sbroffset8_1 = (i[15] & i[14]) & i[0];
	assign simm9_4 = ((((((!i[15] & i[14]) & i[13]) & !i[11]) & !i[10]) & !i[9]) & i[8]) & !i[7];
	assign simm5_0 = ((((!i[14] & !i[13]) & i[11]) & !i[10]) & i[0]) | ((!i[15] & !i[13]) & i[0]);
	assign sjaloffset11_1 = !i[14] & i[13];
	assign sluimm17_12 = ((((((!i[15] & i[14]) & i[13]) & i[7]) | (((!i[15] & i[14]) & i[13]) & !i[8])) | (((!i[15] & i[14]) & i[13]) & i[9])) | (((!i[15] & i[14]) & i[13]) & i[10])) | (((!i[15] & i[14]) & i[13]) & i[11]);
	assign uimm5_0 = ((((i[15] & !i[14]) & !i[13]) & !i[11]) & i[0]) | ((!i[15] & !i[14]) & i[1]);
	assign uswimm6_2 = (i[15] & !i[1]) & !i[0];
	assign uswspimm7_2 = (i[15] & i[14]) & i[1];
	assign o[31] = 1'b0;
	assign o[30] = ((((((i[15] & !i[14]) & !i[13]) & i[10]) & !i[6]) & !i[5]) & i[0]) | (((((i[15] & !i[14]) & !i[13]) & !i[11]) & i[10]) & i[0]);
	assign o[29] = 1'b0;
	assign o[28] = 1'b0;
	assign o[27] = 1'b0;
	assign o[26] = 1'b0;
	assign o[25] = 1'b0;
	assign o[24] = 1'b0;
	assign o[23] = 1'b0;
	assign o[22] = 1'b0;
	assign o[21] = 1'b0;
	assign o[20] = (((((((((((!i[14] & i[12]) & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1];
	assign o[19] = 1'b0;
	assign o[18] = 1'b0;
	assign o[17] = 1'b0;
	assign o[16] = 1'b0;
	assign o[15] = 1'b0;
	assign o[14] = ((((((i[15] & !i[14]) & !i[13]) & !i[11]) & i[0]) | ((((i[15] & !i[14]) & !i[13]) & !i[10]) & i[0])) | ((((i[15] & !i[14]) & !i[13]) & i[6]) & i[0])) | ((((i[15] & !i[14]) & !i[13]) & i[5]) & i[0]);
	assign o[13] = ((((((i[15] & !i[14]) & !i[13]) & i[11]) & !i[10]) & i[0]) | (((((i[15] & !i[14]) & !i[13]) & i[11]) & i[6]) & i[0])) | (i[14] & !i[0]);
	assign o[12] = ((((((((i[15] & !i[14]) & !i[13]) & i[6]) & i[5]) & i[0]) | ((((i[15] & !i[14]) & !i[13]) & !i[11]) & i[0])) | ((((i[15] & !i[14]) & !i[13]) & !i[10]) & i[0])) | ((!i[15] & !i[14]) & i[1])) | ((i[15] & i[14]) & i[13]);
	assign o[11] = 1'b0;
	assign o[10] = 1'b0;
	assign o[9] = 1'b0;
	assign o[8] = 1'b0;
	assign o[7] = 1'b0;
	assign o[6] = ((((((((i[15] & !i[14]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & !i[0]) | (!i[14] & i[13])) | ((i[15] & i[14]) & i[0]);
	assign o[5] = ((((((((i[15] & !i[0]) | ((i[15] & i[11]) & i[10])) | (i[13] & !i[8])) | (i[13] & i[7])) | (i[13] & i[9])) | (i[13] & i[10])) | (i[13] & i[11])) | (!i[14] & i[13])) | (i[15] & i[14]);
	assign o[4] = (((((((((((((!i[14] & !i[11]) & !i[10]) & !i[9]) & !i[8]) & !i[7]) & !i[0]) | ((!i[15] & !i[14]) & !i[0])) | ((!i[14] & i[6]) & !i[0])) | ((!i[15] & i[14]) & i[0])) | ((!i[14] & i[5]) & !i[0])) | ((!i[14] & i[4]) & !i[0])) | ((!i[14] & !i[13]) & i[0])) | ((!i[14] & i[3]) & !i[0])) | ((!i[14] & i[2]) & !i[0]);
	assign o[3] = !i[14] & i[13];
	assign o[2] = ((((((((((((((((((!i[14] & i[12]) & i[11]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1]) | ((((((((!i[14] & i[12]) & i[10]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[9]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[8]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((!i[14] & i[12]) & i[7]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & i[1])) | ((((((((i[15] & !i[14]) & !i[12]) & !i[6]) & !i[5]) & !i[4]) & !i[3]) & !i[2]) & !i[0])) | ((!i[15] & i[13]) & !i[8])) | ((!i[15] & i[13]) & i[7])) | ((!i[15] & i[13]) & i[9])) | ((!i[15] & i[13]) & i[10])) | ((!i[15] & i[13]) & i[11])) | (!i[14] & i[13]);
	assign o[1] = 1'b1;
	assign o[0] = 1'b1;
	assign legal = (((((((((((((((((((((((((((((((((!i[13] & !i[12]) & i[11]) & i[1]) & !i[0]) | ((((!i[13] & !i[12]) & i[6]) & i[1]) & !i[0])) | (((!i[15] & !i[13]) & i[11]) & !i[1])) | ((((!i[13] & !i[12]) & i[5]) & i[1]) & !i[0])) | ((((!i[13] & !i[12]) & i[10]) & i[1]) & !i[0])) | (((!i[15] & !i[13]) & i[6]) & !i[1])) | (((i[15] & !i[12]) & !i[1]) & i[0])) | ((((!i[13] & !i[12]) & i[9]) & i[1]) & !i[0])) | (((!i[12] & i[6]) & !i[1]) & i[0])) | (((!i[15] & !i[13]) & i[5]) & !i[1])) | ((((!i[13] & !i[12]) & i[8]) & i[1]) & !i[0])) | (((!i[12] & i[5]) & !i[1]) & i[0])) | (((!i[15] & !i[13]) & i[10]) & !i[1])) | ((((!i[13] & !i[12]) & i[7]) & i[1]) & !i[0])) | ((((i[12] & i[11]) & !i[10]) & !i[1]) & i[0])) | (((!i[15] & !i[13]) & i[9]) & !i[1])) | ((((!i[13] & !i[12]) & i[4]) & i[1]) & !i[0])) | (((i[13] & i[12]) & !i[1]) & i[0])) | (((!i[15] & !i[13]) & i[8]) & !i[1])) | ((((!i[13] & !i[12]) & i[3]) & i[1]) & !i[0])) | (((i[13] & i[4]) & !i[1]) & i[0])) | ((((!i[13] & !i[12]) & i[2]) & i[1]) & !i[0])) | (((!i[15] & !i[13]) & i[7]) & !i[1])) | (((i[13] & i[3]) & !i[1]) & i[0])) | (((i[13] & i[2]) & !i[1]) & i[0])) | ((i[14] & !i[13]) & !i[1])) | (((!i[14] & !i[12]) & !i[1]) & i[0])) | ((((i[15] & !i[13]) & i[12]) & i[1]) & !i[0])) | ((((!i[15] & !i[13]) & !i[12]) & i[1]) & !i[0])) | (((!i[15] & !i[13]) & i[12]) & !i[1])) | ((i[14] & !i[13]) & !i[0]);
endmodule
module eb1_ifu_iccm_mem (
`ifdef USE_POWER_PINS	
	VPWR,
	VGND,
`endif
	clk,
	active_clk,
	rst_l,
	clk_override,
	iccm_wren,
	iccm_rden,
	iccm_rw_addr,
	iccm_buf_correct_ecc,
	iccm_correction_state,
	iccm_wr_size,
	iccm_wr_data,
	iccm_ext_in_pkt,
	iccm_rd_data,
	iccm_rd_data_ecc,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
`ifdef USE_POWER_PINS
	inout wire VPWR;
	inout wire VGND;
`endif
	input wire clk;
	input wire active_clk;
	input wire rst_l;
	input wire clk_override;
	input wire iccm_wren;
	input wire iccm_rden;
	input wire [pt[936-:9] - 1:1] iccm_rw_addr;
	input wire iccm_buf_correct_ecc;
	input wire iccm_correction_state;
	input wire [2:0] iccm_wr_size;
	input wire [77:0] iccm_wr_data;
	input wire [(pt[909-:9] * 12) - 1:0] iccm_ext_in_pkt;
	output wire [63:0] iccm_rd_data;
	output wire [77:0] iccm_rd_data_ecc;
	input wire scan_mode;
	wire [pt[909-:9] - 1:0] wren_bank;
	wire [pt[909-:9] - 1:0] rden_bank;
	wire [pt[909-:9] - 1:0] iccm_clken;
	wire [((pt[936-:9] - 1) >= pt[945-:9] ? (pt[909-:9] * (((pt[936-:9] - 1) - pt[945-:9]) + 1)) + (pt[945-:9] - 1) : (pt[909-:9] * ((pt[945-:9] - (pt[936-:9] - 1)) + 1)) + (pt[936-:9] - 2)):((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1)] addr_bank;
	wire [(pt[909-:9] * 39) - 1:0] iccm_bank_dout;
	wire [(pt[909-:9] * 39) - 1:0] iccm_bank_dout_fn;
	wire [(pt[909-:9] * 39) - 1:0] iccm_bank_wr_data;
	wire [pt[936-:9] - 1:1] addr_bank_inc;
	wire [pt[954-:9]:2] iccm_rd_addr_hi_q;
	wire [pt[954-:9]:1] iccm_rd_addr_lo_q;
	wire [63:0] iccm_rd_data_pre;
	wire [63:0] iccm_data;
	wire [1:0] addr_incr;
	wire [(pt[909-:9] * 39) - 1:0] iccm_bank_wr_data_vec;
	wire [((pt[936-:9] - 1) >= 2 ? (2 * (pt[936-:9] - 2)) + 1 : (2 * (4 - pt[936-:9])) + (pt[936-:9] - 2)):((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)] redundant_address;
	wire [77:0] redundant_data;
	wire [1:0] redundant_valid;
	wire [pt[909-:9] - 1:0] sel_red1;
	wire [pt[909-:9] - 1:0] sel_red0;
	wire [pt[909-:9] - 1:0] sel_red1_q;
	wire [pt[909-:9] - 1:0] sel_red0_q;
	wire [38:0] redundant_data0_in;
	wire [38:0] redundant_data1_in;
	wire redundant_lru;
	wire redundant_lru_in;
	wire redundant_lru_en;
	wire redundant_data0_en;
	wire redundant_data1_en;
	wire r0_addr_en;
	wire r1_addr_en;
	assign addr_incr[1:0] = (iccm_wr_size[1:0] == 2'b11 ? 2'b10 : 2'b01);
	assign addr_bank_inc[pt[936-:9] - 1:1] = iccm_rw_addr[pt[936-:9] - 1:1] + addr_incr[1:0];
	generate
		genvar i;
		for (i = 0; i < (pt[909-:9] / 2); i = i + 1) begin : mem_bank_data
			assign iccm_bank_wr_data_vec[(2 * i) * 39+:39] = iccm_wr_data[38:0];
			assign iccm_bank_wr_data_vec[((2 * i) + 1) * 39+:39] = iccm_wr_data[77:39];
		end
	endgenerate
	generate
		for (i = 0; i < pt[909-:9]; i = i + 1) begin : mem_bank
			assign wren_bank[i] = iccm_wren & ((iccm_rw_addr[pt[954-:9]:2] == i) | (addr_bank_inc[pt[954-:9]:2] == i));
			assign iccm_bank_wr_data[i * 39+:39] = iccm_bank_wr_data_vec[i * 39+:39];
			assign rden_bank[i] = iccm_rden & ((iccm_rw_addr[pt[954-:9]:2] == i) | (addr_bank_inc[pt[954-:9]:2] == i));
			assign iccm_clken[i] = (wren_bank[i] | rden_bank[i]) | clk_override;
			assign addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) >= pt[945-:9] ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) - 1) : pt[945-:9] - (((pt[936-:9] - 1) >= pt[945-:9] ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) - 1) - (pt[936-:9] - 1))) : (((i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) >= pt[945-:9] ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) - 1) : pt[945-:9] - (((pt[936-:9] - 1) >= pt[945-:9] ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) - 1) - (pt[936-:9] - 1)))) + ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)) - 1)-:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)] = (wren_bank[i] ? iccm_rw_addr[pt[936-:9] - 1:pt[945-:9]] : (addr_bank_inc[pt[954-:9]:2] == i ? addr_bank_inc[pt[936-:9] - 1:pt[945-:9]] : iccm_rw_addr[pt[936-:9] - 1:pt[945-:9]]));
			if (pt[917-:8] == 6) begin : iccm
				ram_64x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 7) begin : iccm
				ram_128x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 8) begin : iccm
				sky130_sram_1kbyte_1rw1r_32x256_8 sram(
					`ifdef USE_POWER_PINS 
					.vccd1(VPWR),
					.vssd1(VGND),
					`endif
					.clk0(clk),
					.csb0(~iccm_clken[i]),
					.web0(~wren_bank[i]),
					.wmask0(4'hf),
					.addr0(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.din0(iccm_bank_wr_data[(i * 39) + 31-:32]),
					.dout0(iccm_bank_dout[(i * 39) + 31-:32]),
					.clk1(clk),
					.csb1(1'b1),
					.addr1(8'h00),
					.dout1()
				);
			end
			else if (pt[917-:8] == 9) begin : iccm
				ram_512x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 10) begin : iccm
				sky130_sram_1kbyte_1rw1r_32x256_8 sram(
					`ifdef USE_POWER_PINS
					.vccd1(VPWR),
					.vssd1(VGND),
					`endif
					.clk0(clk),
					.csb0(~iccm_clken[i]),
					.web0(~wren_bank[i]),
					.wmask0(4'hf),
					.addr0(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.din0(iccm_bank_wr_data[i * 39+:39]),
					.dout0(iccm_bank_dout[i * 39+:39]),
					.clk1(clk),
					.csb1(1'b1),
					.addr1(8'h00),
					.dout1()
				);
			end
			else if (pt[917-:8] == 11) begin : iccm
				ram_2048x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 12) begin : iccm
				ram_4096x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 13) begin : iccm
				ram_8192x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else if (pt[917-:8] == 14) begin : iccm
				ram_16384x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			else begin : iccm
				ram_32768x39 iccm_bank(
					.CLK(clk),
					.ME(iccm_clken[i]),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[936-:9] - 1) >= pt[945-:9] ? pt[945-:9] : pt[936-:9] - 1) + (i * ((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1))+:((pt[936-:9] - 1) >= pt[945-:9] ? ((pt[936-:9] - 1) - pt[945-:9]) + 1 : (pt[945-:9] - (pt[936-:9] - 1)) + 1)]),
					.D(iccm_bank_wr_data[(i * 39) + 38-:39]),
					.Q(iccm_bank_dout[(i * 39) + 38-:39]),
					.ROP(),
					.TEST1(iccm_ext_in_pkt[(i * 12) + 11]),
					.RME(iccm_ext_in_pkt[(i * 12) + 10]),
					.RM(iccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(iccm_ext_in_pkt[(i * 12) + 5]),
					.DS(iccm_ext_in_pkt[(i * 12) + 4]),
					.SD(iccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(iccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(iccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(iccm_ext_in_pkt[i * 12])
				);
			end
			assign sel_red1[i] = redundant_valid[1] & (((iccm_rw_addr[pt[936-:9] - 1:2] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : ((((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1)))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])]) & (iccm_rw_addr[3:2] == i)) | ((addr_bank_inc[pt[936-:9] - 1:2] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : ((((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1)))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])]) & (addr_bank_inc[3:2] == i)));
			assign sel_red0[i] = redundant_valid[0] & (((iccm_rw_addr[pt[936-:9] - 1:2] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : (((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])]) & (iccm_rw_addr[3:2] == i)) | ((addr_bank_inc[pt[936-:9] - 1:2] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : (((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])]) & (addr_bank_inc[3:2] == i)));
			rvdff #(.WIDTH(1)) selred0(
				.rst_l(rst_l),
				.clk(active_clk),
				.din(sel_red0[i]),
				.dout(sel_red0_q[i])
			);
			rvdff #(.WIDTH(1)) selred1(
				.rst_l(rst_l),
				.clk(active_clk),
				.din(sel_red1[i]),
				.dout(sel_red1_q[i])
			);
			assign iccm_bank_dout_fn[(i * 39) + 38-:39] = (({39 {sel_red1_q[i]}} & redundant_data[77-:39]) | ({39 {sel_red0_q[i]}} & redundant_data[38-:39])) | ({39 {~sel_red0_q[i] & ~sel_red1_q[i]}} & iccm_bank_dout[(i * 39) + 38-:39]);
		end
	endgenerate
	assign r0_addr_en = ~redundant_lru & iccm_buf_correct_ecc;
	assign r1_addr_en = redundant_lru & iccm_buf_correct_ecc;
	assign redundant_lru_en = iccm_buf_correct_ecc | (((|sel_red0[pt[909-:9] - 1:0] | |sel_red1[pt[909-:9] - 1:0]) & iccm_rden) & iccm_correction_state);
	assign redundant_lru_in = (iccm_buf_correct_ecc ? ~redundant_lru : (|sel_red0[pt[909-:9] - 1:0] ? 1'b1 : 1'b0));
	rvdffs red_lru(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(redundant_lru_en),
		.din(redundant_lru_in),
		.dout(redundant_lru)
	);
	rvdffs #(.WIDTH(pt[936-:9] - 2)) r0_address(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(r0_addr_en),
		.din(iccm_rw_addr[pt[936-:9] - 1:2]),
		.dout(redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : (((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])])
	);
	rvdffs #(.WIDTH(pt[936-:9] - 2)) r1_address(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(r1_addr_en),
		.din(iccm_rw_addr[pt[936-:9] - 1:2]),
		.dout(redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : ((((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1) - (pt[936-:9] - 1)))) + ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9])])
	);
	rvdffs #(.WIDTH(1)) r0_valid(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(r0_addr_en),
		.din(1'b1),
		.dout(redundant_valid[0])
	);
	rvdffs #(.WIDTH(1)) r1_valid(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(r1_addr_en),
		.din(1'b1),
		.dout(redundant_valid[1])
	);
	assign redundant_data0_en = ((((iccm_rw_addr[pt[936-:9] - 1:3] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : (((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])]) & ((iccm_rw_addr[2] == redundant_address[((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)]) | (iccm_wr_size[1:0] == 2'b11))) & redundant_valid[0]) & iccm_wren) | (~redundant_lru & iccm_buf_correct_ecc);
	assign redundant_data0_in[38:0] = (((iccm_rw_addr[2] == redundant_address[((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)]) & iccm_rw_addr[2]) | (redundant_address[((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)] & (iccm_wr_size[1:0] == 2'b11)) ? iccm_wr_data[77:39] : iccm_wr_data[38:0]);
	rvdffs #(.WIDTH(39)) r0_data(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(redundant_data0_en),
		.din(redundant_data0_in[38:0]),
		.dout(redundant_data[38-:39])
	);
	assign redundant_data1_en = ((((iccm_rw_addr[pt[936-:9] - 1:3] == redundant_address[((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) - (pt[936-:9] - 1))) : ((((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) : 2 - (((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 1 : ((pt[936-:9] - 1) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1) - (pt[936-:9] - 1)))) + ((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])) - 1)-:((pt[936-:9] - 1) >= 3 ? pt[936-:9] - 3 : 5 - pt[936-:9])]) & ((iccm_rw_addr[2] == redundant_address[((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)]) | (iccm_wr_size[1:0] == 2'b11))) & redundant_valid[1]) & iccm_wren) | (redundant_lru & iccm_buf_correct_ecc);
	assign redundant_data1_in[38:0] = (((iccm_rw_addr[2] == redundant_address[((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)]) & iccm_rw_addr[2]) | (redundant_address[((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) + ((pt[936-:9] - 1) >= 2 ? 2 : pt[936-:9] - 1)] & (iccm_wr_size[1:0] == 2'b11)) ? iccm_wr_data[77:39] : iccm_wr_data[38:0]);
	rvdffs #(.WIDTH(39)) r1_data(
		.rst_l(rst_l),
		.clk(active_clk),
		.en(redundant_data1_en),
		.din(redundant_data1_in[38:0]),
		.dout(redundant_data[77-:39])
	);
	rvdffs #(.WIDTH(pt[954-:9])) rd_addr_lo_ff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din(iccm_rw_addr[pt[954-:9]:1]),
		.dout(iccm_rd_addr_lo_q[pt[954-:9]:1]),
		.en(1'b1)
	);
	rvdffs #(.WIDTH(pt[961-:7])) rd_addr_hi_ff(
		.rst_l(rst_l),
		.clk(active_clk),
		.din(addr_bank_inc[pt[954-:9]:2]),
		.dout(iccm_rd_addr_hi_q[pt[954-:9]:2]),
		.en(1'b1)
	);
	assign iccm_rd_data_pre[63:0] = {iccm_bank_dout_fn[(iccm_rd_addr_hi_q * 39) + 31-:32], iccm_bank_dout_fn[(iccm_rd_addr_lo_q[pt[954-:9]:2] * 39) + 31-:32]};
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	assign iccm_data[63:0] = sv2v_cast_64({16'b0000000000000000, iccm_rd_data_pre[63:0] >> (16 * iccm_rd_addr_lo_q[1])});
	assign iccm_rd_data[63:0] = {iccm_data[63:0]};
	assign iccm_rd_data_ecc[77:0] = {iccm_bank_dout_fn[(iccm_rd_addr_hi_q * 39) + 38-:39], iccm_bank_dout_fn[(iccm_rd_addr_lo_q[pt[954-:9]:2] * 39) + 38-:39]};
endmodule
module eb1_ifu_ifc_ctl (
	clk,
	free_l2clk,
	rst_l,
	scan_mode,
	ic_hit_f,
	ifu_ic_mb_empty,
	ifu_fb_consume1,
	ifu_fb_consume2,
	dec_tlu_flush_noredir_wb,
	exu_flush_final,
	exu_flush_path_final,
	ifu_bp_hit_taken_f,
	ifu_bp_btb_target_f,
	ic_dma_active,
	ic_write_stall,
	dma_iccm_stall_any,
	dec_tlu_mrac_ff,
	ifc_fetch_addr_f,
	ifc_fetch_addr_bf,
	ifc_fetch_req_f,
	ifu_pmu_fetch_stall,
	ifc_fetch_uncacheable_bf,
	ifc_fetch_req_bf,
	ifc_fetch_req_bf_raw,
	ifc_iccm_access_bf,
	ifc_region_acc_fault_bf,
	ifc_dma_access_ok
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire free_l2clk;
	input wire rst_l;
	input wire scan_mode;
	input wire ic_hit_f;
	input wire ifu_ic_mb_empty;
	input wire ifu_fb_consume1;
	input wire ifu_fb_consume2;
	input wire dec_tlu_flush_noredir_wb;
	input wire exu_flush_final;
	input wire [31:1] exu_flush_path_final;
	input wire ifu_bp_hit_taken_f;
	input wire [31:1] ifu_bp_btb_target_f;
	input wire ic_dma_active;
	input wire ic_write_stall;
	input wire dma_iccm_stall_any;
	input wire [31:0] dec_tlu_mrac_ff;
	output wire [31:1] ifc_fetch_addr_f;
	output wire [31:1] ifc_fetch_addr_bf;
	output wire ifc_fetch_req_f;
	output wire ifu_pmu_fetch_stall;
	output wire ifc_fetch_uncacheable_bf;
	output wire ifc_fetch_req_bf;
	output wire ifc_fetch_req_bf_raw;
	output wire ifc_iccm_access_bf;
	output wire ifc_region_acc_fault_bf;
	output wire ifc_dma_access_ok;
	wire [31:1] fetch_addr_bf;
	wire [31:1] fetch_addr_next;
	wire [3:0] fb_write_f;
	wire [3:0] fb_write_ns;
	wire fb_full_f_ns;
	wire fb_full_f;
	wire fb_right;
	wire fb_right2;
	wire fb_left;
	wire wfm;
	wire idle;
	wire sel_last_addr_bf;
	wire sel_next_addr_bf;
	wire miss_f;
	wire miss_a;
	wire flush_fb;
	wire dma_iccm_stall_any_f;
	wire mb_empty_mod;
	wire goto_idle;
	wire leave_idle;
	wire fetch_bf_en;
	wire line_wrap;
	wire fetch_addr_next_1;
	wire [1:0] state;
	wire [1:0] next_state;
	wire dma_stall;
	assign dma_stall = ic_dma_active | dma_iccm_stall_any_f;
	generate
		if (pt[2130-:5] == 1) begin
			wire sel_btb_addr_bf;
			assign sel_last_addr_bf = ~exu_flush_final & (~ifc_fetch_req_f | ~ic_hit_f);
			assign sel_btb_addr_bf = ((~exu_flush_final & ifc_fetch_req_f) & ifu_bp_hit_taken_f) & ic_hit_f;
			assign sel_next_addr_bf = ((~exu_flush_final & ifc_fetch_req_f) & ~ifu_bp_hit_taken_f) & ic_hit_f;
			assign fetch_addr_bf[31:1] = ((({31 {exu_flush_final}} & exu_flush_path_final[31:1]) | ({31 {sel_last_addr_bf}} & ifc_fetch_addr_f[31:1])) | ({31 {sel_btb_addr_bf}} & {ifu_bp_btb_target_f[31:1]})) | ({31 {sel_next_addr_bf}} & {fetch_addr_next[31:1]});
		end
		else begin
			assign sel_last_addr_bf = ~exu_flush_final & (~ifc_fetch_req_f | ~ic_hit_f);
			assign sel_next_addr_bf = (~exu_flush_final & ifc_fetch_req_f) & ic_hit_f;
			assign fetch_addr_bf[31:1] = (({31 {exu_flush_final}} & exu_flush_path_final[31:1]) | ({31 {sel_last_addr_bf}} & ifc_fetch_addr_f[31:1])) | ({31 {sel_next_addr_bf}} & {fetch_addr_next[31:1]});
		end
	endgenerate
	assign fetch_addr_next[31:1] = {{ifc_fetch_addr_f[31:2]} + 31'b0000000000000000000000000000001, fetch_addr_next_1};
	assign line_wrap = fetch_addr_next[pt[998-:7]] ^ ifc_fetch_addr_f[pt[998-:7]];
	assign fetch_addr_next_1 = (line_wrap ? 1'b0 : ifc_fetch_addr_f[1]);
	assign ifc_fetch_req_bf_raw = ~idle;
	assign ifc_fetch_req_bf = (((ifc_fetch_req_bf_raw & ~(fb_full_f_ns & ~(ifu_fb_consume2 | ifu_fb_consume1))) & ~dma_stall) & ~ic_write_stall) & ~dec_tlu_flush_noredir_wb;
	assign fetch_bf_en = exu_flush_final | ifc_fetch_req_f;
	assign miss_f = (ifc_fetch_req_f & ~ic_hit_f) & ~exu_flush_final;
	assign mb_empty_mod = (((ifu_ic_mb_empty | exu_flush_final) & ~dma_stall) & ~miss_f) & ~miss_a;
	assign goto_idle = exu_flush_final & dec_tlu_flush_noredir_wb;
	assign leave_idle = (exu_flush_final & ~dec_tlu_flush_noredir_wb) & idle;
	assign next_state[1] = (((~state[1] & state[0]) & miss_f) & ~goto_idle) | ((state[1] & ~mb_empty_mod) & ~goto_idle);
	assign next_state[0] = (~goto_idle & leave_idle) | (state[0] & ~goto_idle);
	assign flush_fb = exu_flush_final;
	assign fb_right = ((ifu_fb_consume1 & ~ifu_fb_consume2) & (~ifc_fetch_req_f | miss_f)) | (ifu_fb_consume2 & ifc_fetch_req_f);
	assign fb_right2 = ifu_fb_consume2 & (~ifc_fetch_req_f | miss_f);
	assign fb_left = (ifc_fetch_req_f & ~(ifu_fb_consume1 | ifu_fb_consume2)) & ~miss_f;
	assign fb_write_ns[3:0] = (((({4 {flush_fb}} & 4'b0001) | ({4 {~flush_fb & fb_right}} & {1'b0, fb_write_f[3:1]})) | ({4 {~flush_fb & fb_right2}} & {2'b00, fb_write_f[3:2]})) | ({4 {~flush_fb & fb_left}} & {fb_write_f[2:0], 1'b0})) | ({4 {((~flush_fb & ~fb_right) & ~fb_right2) & ~fb_left}} & fb_write_f[3:0]);
	assign fb_full_f_ns = fb_write_ns[3];
	localparam [1:0] IDLE = 2'b00;
	assign idle = state == IDLE;
	localparam [1:0] WFM = 2'b11;
	assign wfm = state == WFM;
	rvdffie #(.WIDTH(10)) fbwrite_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({dma_iccm_stall_any, miss_f, ifc_fetch_req_bf, next_state[1:0], fb_full_f_ns, fb_write_ns[3:0]}),
		.dout({dma_iccm_stall_any_f, miss_a, ifc_fetch_req_f, state[1:0], fb_full_f, fb_write_f[3:0]})
	);
	assign ifu_pmu_fetch_stall = wfm | (ifc_fetch_req_bf_raw & ((fb_full_f & ~((ifu_fb_consume2 | ifu_fb_consume1) | exu_flush_final)) | dma_stall));
	assign ifc_fetch_addr_bf[31:1] = fetch_addr_bf[31:1];
	rvdffpcie #(.WIDTH(31)) faddrf1_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(fetch_bf_en),
		.din(fetch_addr_bf[31:1]),
		.dout(ifc_fetch_addr_f[31:1])
	);
	generate
		if (pt[927-:5]) begin
			wire iccm_acc_in_region_bf;
			wire iccm_acc_in_range_bf;
			rvrangecheck #(
				.CCM_SADR(pt[887-:36]),
				.CCM_SIZE(pt[851-:14])
			) iccm_rangecheck(
				.addr({ifc_fetch_addr_bf[31:1], 1'b0}),
				.in_range(iccm_acc_in_range_bf),
				.in_region(iccm_acc_in_region_bf)
			);
			assign ifc_iccm_access_bf = iccm_acc_in_range_bf;
			assign ifc_dma_access_ok = ((((~ifc_iccm_access_bf | (fb_full_f & ~(ifu_fb_consume2 | ifu_fb_consume1))) | (wfm & ~ifc_fetch_req_bf)) | idle) & ~exu_flush_final) | dma_iccm_stall_any_f;
			assign ifc_region_acc_fault_bf = ~iccm_acc_in_range_bf & iccm_acc_in_region_bf;
		end
		else begin
			assign ifc_iccm_access_bf = 1'b0;
			assign ifc_dma_access_ok = 1'b0;
			assign ifc_region_acc_fault_bf = 1'b0;
		end
	endgenerate
	assign ifc_fetch_uncacheable_bf = ~dec_tlu_mrac_ff[{ifc_fetch_addr_bf[31:28], 1'b0}];
endmodule
module eb1_ifu_mem_ctl (
	clk,
	active_clk,
	free_l2clk,
	rst_l,
	exu_flush_final,
	dec_tlu_flush_lower_wb,
	dec_tlu_flush_err_wb,
	dec_tlu_i0_commit_cmt,
	dec_tlu_force_halt,
	ifc_fetch_addr_bf,
	ifc_fetch_uncacheable_bf,
	ifc_fetch_req_bf,
	ifc_fetch_req_bf_raw,
	ifc_iccm_access_bf,
	ifc_region_acc_fault_bf,
	ifc_dma_access_ok,
	dec_tlu_fence_i_wb,
	ifu_bp_hit_taken_f,
	ifu_bp_inst_mask_f,
	ifu_miss_state_idle,
	ifu_ic_mb_empty,
	ic_dma_active,
	ic_write_stall,
	ifu_pmu_ic_miss,
	ifu_pmu_ic_hit,
	ifu_pmu_bus_error,
	ifu_pmu_bus_busy,
	ifu_pmu_bus_trxn,
	ifu_axi_awvalid,
	ifu_axi_awid,
	ifu_axi_awaddr,
	ifu_axi_awregion,
	ifu_axi_awlen,
	ifu_axi_awsize,
	ifu_axi_awburst,
	ifu_axi_awlock,
	ifu_axi_awcache,
	ifu_axi_awprot,
	ifu_axi_awqos,
	ifu_axi_wvalid,
	ifu_axi_wdata,
	ifu_axi_wstrb,
	ifu_axi_wlast,
	ifu_axi_bready,
	ifu_axi_arvalid,
	ifu_axi_arready,
	ifu_axi_arid,
	ifu_axi_araddr,
	ifu_axi_arregion,
	ifu_axi_arlen,
	ifu_axi_arsize,
	ifu_axi_arburst,
	ifu_axi_arlock,
	ifu_axi_arcache,
	ifu_axi_arprot,
	ifu_axi_arqos,
	ifu_axi_rvalid,
	ifu_axi_rready,
	ifu_axi_rid,
	ifu_axi_rdata,
	ifu_axi_rresp,
	ifu_bus_clk_en,
	dma_iccm_req,
	dma_mem_addr,
	dma_mem_sz,
	dma_mem_write,
	dma_mem_wdata,
	dma_mem_tag,
	iccm_dma_ecc_error,
	iccm_dma_rvalid,
	iccm_dma_rdata,
	iccm_dma_rtag,
	iccm_ready,
	ic_rw_addr,
	ic_wr_en,
	ic_rd_en,
	ic_wr_data,
	ic_rd_data,
	ic_debug_rd_data,
	ictag_debug_rd_data,
	ic_debug_wr_data,
	ifu_ic_debug_rd_data,
	ic_eccerr,
	ic_parerr,
	ic_debug_addr,
	ic_debug_rd_en,
	ic_debug_wr_en,
	ic_debug_tag_array,
	ic_debug_way,
	ic_tag_valid,
	ic_rd_hit,
	ic_tag_perr,
	iccm_rw_addr,
	iccm_wren,
	iccm_rden,
	iccm_wr_data,
	iccm_wr_size,
	iccm_rd_data,
	iccm_rd_data_ecc,
	ifu_fetch_val,
	ic_hit_f,
	ic_access_fault_f,
	ic_access_fault_type_f,
	iccm_rd_ecc_single_err,
	iccm_rd_ecc_double_err,
	ic_error_start,
	ifu_async_error_start,
	iccm_dma_sb_error,
	ic_fetch_val_f,
	ic_data_f,
	ic_premux_data,
	ic_sel_premux_data,
	dec_tlu_ic_diag_pkt,
	dec_tlu_core_ecc_disable,
	ifu_ic_debug_rd_data_valid,
	iccm_buf_correct_ecc,
	iccm_correction_state,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire active_clk;
	input wire free_l2clk;
	input wire rst_l;
	input wire exu_flush_final;
	input wire dec_tlu_flush_lower_wb;
	input wire dec_tlu_flush_err_wb;
	input wire dec_tlu_i0_commit_cmt;
	input wire dec_tlu_force_halt;
	input wire [31:1] ifc_fetch_addr_bf;
	input wire ifc_fetch_uncacheable_bf;
	input wire ifc_fetch_req_bf;
	input wire ifc_fetch_req_bf_raw;
	input wire ifc_iccm_access_bf;
	input wire ifc_region_acc_fault_bf;
	input wire ifc_dma_access_ok;
	input wire dec_tlu_fence_i_wb;
	input wire ifu_bp_hit_taken_f;
	input wire ifu_bp_inst_mask_f;
	output wire ifu_miss_state_idle;
	output wire ifu_ic_mb_empty;
	output wire ic_dma_active;
	output wire ic_write_stall;
	output wire ifu_pmu_ic_miss;
	output wire ifu_pmu_ic_hit;
	output wire ifu_pmu_bus_error;
	output wire ifu_pmu_bus_busy;
	output wire ifu_pmu_bus_trxn;
	output wire ifu_axi_awvalid;
	output wire [pt[826-:8] - 1:0] ifu_axi_awid;
	output wire [31:0] ifu_axi_awaddr;
	output wire [3:0] ifu_axi_awregion;
	output wire [7:0] ifu_axi_awlen;
	output wire [2:0] ifu_axi_awsize;
	output wire [1:0] ifu_axi_awburst;
	output wire ifu_axi_awlock;
	output wire [3:0] ifu_axi_awcache;
	output wire [2:0] ifu_axi_awprot;
	output wire [3:0] ifu_axi_awqos;
	output wire ifu_axi_wvalid;
	output wire [63:0] ifu_axi_wdata;
	output wire [7:0] ifu_axi_wstrb;
	output wire ifu_axi_wlast;
	output wire ifu_axi_bready;
	output wire ifu_axi_arvalid;
	input wire ifu_axi_arready;
	output wire [pt[826-:8] - 1:0] ifu_axi_arid;
	output wire [31:0] ifu_axi_araddr;
	output wire [3:0] ifu_axi_arregion;
	output wire [7:0] ifu_axi_arlen;
	output wire [2:0] ifu_axi_arsize;
	output wire [1:0] ifu_axi_arburst;
	output wire ifu_axi_arlock;
	output wire [3:0] ifu_axi_arcache;
	output wire [2:0] ifu_axi_arprot;
	output wire [3:0] ifu_axi_arqos;
	input wire ifu_axi_rvalid;
	output wire ifu_axi_rready;
	input wire [pt[826-:8] - 1:0] ifu_axi_rid;
	input wire [63:0] ifu_axi_rdata;
	input wire [1:0] ifu_axi_rresp;
	input wire ifu_bus_clk_en;
	input wire dma_iccm_req;
	input wire [31:0] dma_mem_addr;
	input wire [2:0] dma_mem_sz;
	input wire dma_mem_write;
	input wire [63:0] dma_mem_wdata;
	input wire [2:0] dma_mem_tag;
	output wire iccm_dma_ecc_error;
	output wire iccm_dma_rvalid;
	output wire [63:0] iccm_dma_rdata;
	output wire [2:0] iccm_dma_rtag;
	output wire iccm_ready;
	output wire [31:1] ic_rw_addr;
	output wire [pt[1060-:7] - 1:0] ic_wr_en;
	output wire ic_rd_en;
	output wire [(pt[1189-:7] * 71) - 1:0] ic_wr_data;
	input wire [63:0] ic_rd_data;
	input wire [70:0] ic_debug_rd_data;
	input wire [25:0] ictag_debug_rd_data;
	output wire [70:0] ic_debug_wr_data;
	output wire [70:0] ifu_ic_debug_rd_data;
	input wire [pt[1189-:7] - 1:0] ic_eccerr;
	input wire [pt[1189-:7] - 1:0] ic_parerr;
	output wire [pt[1104-:9]:3] ic_debug_addr;
	output wire ic_debug_rd_en;
	output wire ic_debug_wr_en;
	output wire ic_debug_tag_array;
	output wire [pt[1060-:7] - 1:0] ic_debug_way;
	output wire [pt[1060-:7] - 1:0] ic_tag_valid;
	input wire [pt[1060-:7] - 1:0] ic_rd_hit;
	input wire ic_tag_perr;
	output wire [pt[936-:9] - 1:1] iccm_rw_addr;
	output wire iccm_wren;
	output wire iccm_rden;
	output wire [77:0] iccm_wr_data;
	output wire [2:0] iccm_wr_size;
	input wire [63:0] iccm_rd_data;
	input wire [77:0] iccm_rd_data_ecc;
	input wire [1:0] ifu_fetch_val;
	output wire ic_hit_f;
	output wire [1:0] ic_access_fault_f;
	output wire [1:0] ic_access_fault_type_f;
	output wire iccm_rd_ecc_single_err;
	output wire [1:0] iccm_rd_ecc_double_err;
	output wire ic_error_start;
	output wire ifu_async_error_start;
	output wire iccm_dma_sb_error;
	output wire [1:0] ic_fetch_val_f;
	output wire [31:0] ic_data_f;
	output wire [63:0] ic_premux_data;
	output wire ic_sel_premux_data;
	input wire [89:0] dec_tlu_ic_diag_pkt;
	input wire dec_tlu_core_ecc_disable;
	output wire ifu_ic_debug_rd_data_valid;
	output wire iccm_buf_correct_ecc;
	output reg iccm_correction_state;
	input wire scan_mode;
	localparam NUM_OF_BEATS = 8;
	wire [31:3] ifu_ic_req_addr_f;
	wire uncacheable_miss_in;
	wire uncacheable_miss_ff;
	wire bus_ifu_wr_en;
	wire bus_ifu_wr_en_ff;
	wire bus_ifu_wr_en_ff_q;
	wire bus_ifu_wr_en_ff_wo_err;
	wire [pt[1060-:7] - 1:0] bus_ic_wr_en;
	wire reset_tag_valid_for_miss;
	reg [pt[1027-:7] - 1:0] way_status;
	wire [pt[1027-:7] - 1:0] way_status_mb_in;
	wire [pt[1027-:7] - 1:0] way_status_rep_new;
	wire [pt[1027-:7] - 1:0] way_status_mb_ff;
	wire [pt[1027-:7] - 1:0] way_status_new;
	wire [pt[1027-:7] - 1:0] way_status_hit_new;
	wire [pt[1027-:7] - 1:0] way_status_new_w_debug;
	wire [pt[1060-:7] - 1:0] tagv_mb_in;
	wire [pt[1060-:7] - 1:0] tagv_mb_ff;
	wire ifu_wr_data_comb_err;
	wire ifu_byp_data_err_new;
	wire [1:0] ifu_byp_data_err_f;
	wire ifu_wr_cumulative_err_data;
	wire ifu_wr_cumulative_err;
	wire ifu_wr_data_comb_err_ff;
	wire scnd_miss_index_match;
	wire ifc_dma_access_q_ok;
	wire ifc_iccm_access_f;
	wire ifc_region_acc_fault_f;
	wire ifc_region_acc_fault_final_f;
	wire [1:0] ifc_bus_acc_fault_f;
	wire ic_act_miss_f;
	wire ic_miss_under_miss_f;
	wire ic_ignore_2nd_miss_f;
	wire ic_act_hit_f;
	wire miss_pending;
	wire [31:1] imb_in;
	wire [31:1] imb_ff;
	wire [31:pt[1182-:8] + 1] miss_addr_in;
	wire [31:pt[1182-:8] + 1] miss_addr;
	wire miss_wrap_f;
	wire flush_final_f;
	wire ifc_fetch_req_f;
	wire ifc_fetch_req_f_raw;
	wire fetch_req_f_qual;
	wire ifc_fetch_req_qual_bf;
	wire [pt[1060-:7] - 1:0] replace_way_mb_any;
	wire last_beat;
	wire reset_beat_cnt;
	wire [pt[1182-:8]:3] ic_req_addr_bits_hi_3;
	wire [pt[1182-:8]:3] ic_wr_addr_bits_hi_3;
	wire [31:1] ifu_fetch_addr_int_f;
	wire [31:1] ifu_ic_rw_int_addr;
	wire crit_wd_byp_ok_ff;
	wire ic_crit_wd_rdy_new_ff;
	wire [79:0] ic_byp_data_only_pre_new;
	wire [79:0] ic_byp_data_only_new;
	wire ic_byp_hit_f;
	wire ic_valid;
	wire ic_valid_ff;
	wire reset_all_tags;
	wire ic_valid_w_debug;
	wire [pt[1060-:7] - 1:0] ifu_tag_wren;
	wire [pt[1060-:7] - 1:0] ifu_tag_wren_ff;
	wire [pt[1060-:7] - 1:0] ic_debug_tag_wr_en;
	wire [pt[1060-:7] - 1:0] ifu_tag_wren_w_debug;
	wire [pt[1060-:7] - 1:0] ic_debug_way_ff;
	wire ic_debug_rd_en_ff;
	wire fetch_bf_f_c1_clken;
	wire fetch_bf_f_c1_clk;
	wire debug_c1_clken;
	wire debug_c1_clk;
	wire reset_ic_in;
	wire reset_ic_ff;
	wire [pt[1182-:8]:1] vaddr_f;
	wire [31:1] ifu_status_wr_addr;
	wire sel_mb_addr;
	wire sel_mb_addr_ff;
	wire sel_mb_status_addr;
	wire [63:0] ic_final_data;
	wire [pt[1104-:9]:pt[998-:7]] ifu_ic_rw_int_addr_ff;
	wire [pt[1104-:9]:pt[998-:7]] ifu_status_wr_addr_ff;
	wire [pt[1104-:9]:pt[998-:7]] ifu_ic_rw_int_addr_w_debug;
	wire [pt[1104-:9]:pt[998-:7]] ifu_status_wr_addr_w_debug;
	wire [pt[1027-:7] - 1:0] way_status_new_ff;
	wire way_status_wr_en_ff;
	wire [(pt[1015-:17] * pt[1027-:7]) - 1:0] way_status_out;
	wire [1:0] ic_debug_way_enc;
	wire [pt[826-:8] - 1:0] ifu_bus_rid_ff;
	wire fetch_req_icache_f;
	wire fetch_req_iccm_f;
	wire ic_iccm_hit_f;
	wire fetch_uncacheable_ff;
	wire way_status_wr_en;
	wire sel_byp_data;
	wire sel_ic_data;
	wire sel_iccm_data;
	wire ic_rd_parity_final_err;
	wire ic_act_miss_f_delayed;
	wire bus_ifu_wr_data_error;
	wire bus_ifu_wr_data_error_ff;
	wire way_status_wr_en_w_debug;
	wire ic_debug_tag_val_rd_out;
	wire ifu_pmu_ic_miss_in;
	wire ifu_pmu_ic_hit_in;
	wire ifu_pmu_bus_error_in;
	wire ifu_pmu_bus_trxn_in;
	wire ifu_pmu_bus_busy_in;
	wire ic_debug_ict_array_sel_in;
	wire ic_debug_ict_array_sel_ff;
	wire debug_data_clken;
	wire last_data_recieved_in;
	wire last_data_recieved_ff;
	wire ifu_bus_rvalid;
	wire ifu_bus_rvalid_ff;
	wire ifu_bus_rvalid_unq_ff;
	wire ifu_bus_arready_unq;
	wire ifu_bus_arready_unq_ff;
	wire ifu_bus_arvalid;
	wire ifu_bus_arvalid_ff;
	wire ifu_bus_arready;
	wire ifu_bus_arready_ff;
	wire [63:0] ifu_bus_rdata_ff;
	wire [1:0] ifu_bus_rresp_ff;
	wire ifu_bus_rsp_valid;
	wire ifu_bus_rsp_ready;
	wire [pt[826-:8] - 1:0] ifu_bus_rsp_tag;
	wire [63:0] ifu_bus_rsp_rdata;
	wire [1:0] ifu_bus_rsp_opc;
	wire [pt[1084-:8] - 1:0] write_fill_data;
	wire [pt[1084-:8] - 1:0] wr_data_c1_clk;
	wire [pt[1084-:8] - 1:0] ic_miss_buff_data_valid_in;
	wire [pt[1084-:8] - 1:0] ic_miss_buff_data_valid;
	wire [pt[1084-:8] - 1:0] ic_miss_buff_data_error_in;
	wire [pt[1084-:8] - 1:0] ic_miss_buff_data_error;
	wire [pt[1182-:8]:1] byp_fetch_index;
	wire [pt[1182-:8]:2] byp_fetch_index_0;
	wire [pt[1182-:8]:2] byp_fetch_index_1;
	wire [pt[1182-:8]:3] byp_fetch_index_inc;
	wire [pt[1182-:8]:2] byp_fetch_index_inc_0;
	wire [pt[1182-:8]:2] byp_fetch_index_inc_1;
	wire miss_buff_hit_unq_f;
	wire stream_hit_f;
	wire stream_miss_f;
	wire stream_eol_f;
	wire crit_byp_hit_f;
	wire [pt[826-:8] - 1:0] other_tag;
	wire [((2 * pt[1084-:8]) * 32) - 1:0] ic_miss_buff_data;
	wire [63:0] ic_miss_buff_half;
	wire scnd_miss_req;
	wire scnd_miss_req_q;
	wire scnd_miss_req_in;
	wire [pt[936-:9] - 1:2] iccm_ecc_corr_index_ff;
	wire [pt[936-:9] - 1:2] iccm_ecc_corr_index_in;
	wire [38:0] iccm_ecc_corr_data_ff;
	wire iccm_ecc_write_status;
	wire iccm_rd_ecc_single_err_ff;
	wire iccm_error_start;
	reg perr_state_en;
	reg miss_state_en;
	wire busclk;
	wire busclk_force;
	wire busclk_reset;
	wire bus_ifu_bus_clk_en_ff;
	wire bus_ifu_bus_clk_en;
	wire ifc_bus_ic_req_ff_in;
	wire ifu_bus_cmd_valid;
	wire ifu_bus_cmd_ready;
	wire bus_inc_data_beat_cnt;
	wire bus_reset_data_beat_cnt;
	wire bus_hold_data_beat_cnt;
	wire bus_inc_cmd_beat_cnt;
	wire bus_reset_cmd_beat_cnt_0;
	wire bus_reset_cmd_beat_cnt_secondlast;
	wire bus_hold_cmd_beat_cnt;
	wire [pt[1174-:8] - 1:0] bus_new_data_beat_count;
	wire [pt[1174-:8] - 1:0] bus_data_beat_count;
	wire [pt[1174-:8] - 1:0] bus_new_cmd_beat_count;
	wire [pt[1174-:8] - 1:0] bus_cmd_beat_count;
	wire [pt[1174-:8] - 1:0] bus_new_rd_addr_count;
	wire [pt[1174-:8] - 1:0] bus_rd_addr_count;
	wire bus_cmd_sent;
	wire bus_last_data_beat;
	wire [pt[1060-:7] - 1:0] bus_wren;
	wire [pt[1060-:7] - 1:0] bus_wren_last;
	wire [pt[1060-:7] - 1:0] wren_reset_miss;
	wire ifc_dma_access_ok_d;
	wire ifc_dma_access_ok_prev;
	wire bus_cmd_req_in;
	wire bus_cmd_req_hold;
	wire second_half_available;
	wire write_ic_16_bytes;
	wire ifc_region_acc_fault_final_bf;
	wire ifc_region_acc_fault_memory_bf;
	wire ifc_region_acc_fault_memory_f;
	wire ifc_region_acc_okay;
	wire iccm_correct_ecc;
	wire dma_sb_err_state;
	wire dma_sb_err_state_ff;
	wire two_byte_instr;
	wire [2:0] miss_state;
	reg [2:0] miss_nxtstate;
	wire [1:0] err_stop_state;
	reg [1:0] err_stop_nxtstate;
	reg err_stop_state_en;
	reg err_stop_fetch;
	wire ic_crit_wd_rdy;
	wire ifu_bp_hit_taken_q_f;
	wire ifu_bus_rvalid_unq;
	wire bus_cmd_beat_en;
	assign fetch_bf_f_c1_clken = (((ifc_fetch_req_bf_raw | ifc_fetch_req_f) | miss_pending) | exu_flush_final) | scnd_miss_req;
	assign debug_c1_clken = ic_debug_rd_en | ic_debug_wr_en;
	rvclkhdr fetch_bf_f_c1_cgc(
		.en(fetch_bf_f_c1_clken),
		.l1clk(fetch_bf_f_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr debug_c1_cgc(
		.en(debug_c1_clken),
		.l1clk(debug_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	wire [1:0] iccm_single_ecc_error;
	wire dma_iccm_req_f;
	assign iccm_dma_sb_error = |iccm_single_ecc_error[1:0] & dma_iccm_req_f;
	assign ifu_async_error_start = iccm_rd_ecc_single_err | ic_error_start;
	wire [2:0] perr_state;
	reg [2:0] perr_nxtstate;
	localparam [2:0] DMA_SB_ERR = 3'b100;
	localparam [1:0] ERR_STOP_FETCH = 2'b11;
	assign ic_dma_active = (((iccm_correct_ecc | (perr_state == DMA_SB_ERR)) | (err_stop_state == ERR_STOP_FETCH)) | err_stop_fetch) | dec_tlu_flush_err_wb;
	localparam [2:0] SCND_MISS = 3'b101;
	assign scnd_miss_req_in = (((((ifu_bus_rsp_valid & bus_ifu_bus_clk_en) & ifu_bus_rsp_ready) & &bus_new_data_beat_count[pt[1174-:8] - 1:0]) & ~uncacheable_miss_ff) & ((miss_state == SCND_MISS) | (miss_nxtstate == SCND_MISS))) & ~exu_flush_final;
	assign ifu_bp_hit_taken_q_f = ifu_bp_hit_taken_f & ic_hit_f;
	localparam [2:0] CRIT_BYP_OK = 3'b001;
	localparam [2:0] CRIT_WRD_RDY = 3'b100;
	localparam [2:0] HIT_U_MISS = 3'b010;
	localparam [2:0] IDLE = 3'b000;
	localparam [2:0] MISS_WAIT = 3'b011;
	localparam [2:0] STALL_SCND_MISS = 3'b111;
	localparam [2:0] STREAM = 3'b110;
	always @(*) begin : MISS_SM
		miss_nxtstate = IDLE;
		miss_state_en = 1'b0;
		case (miss_state)
			IDLE: begin : idle
				miss_nxtstate = (ic_act_miss_f & ~exu_flush_final ? CRIT_BYP_OK : HIT_U_MISS);
				miss_state_en = ic_act_miss_f & ~dec_tlu_force_halt;
			end
			CRIT_BYP_OK: begin : crit_byp_ok
				miss_nxtstate = (dec_tlu_force_halt ? IDLE : ((ic_byp_hit_f & (last_data_recieved_ff | (bus_ifu_wr_en_ff & last_beat))) & uncacheable_miss_ff ? IDLE : ((ic_byp_hit_f & ~last_data_recieved_ff) & uncacheable_miss_ff ? MISS_WAIT : (((~ic_byp_hit_f & ~exu_flush_final) & (bus_ifu_wr_en_ff & last_beat)) & uncacheable_miss_ff ? CRIT_WRD_RDY : ((bus_ifu_wr_en_ff & last_beat) & ~uncacheable_miss_ff ? IDLE : ((((ic_byp_hit_f & ~exu_flush_final) & ~(bus_ifu_wr_en_ff & last_beat)) & ~ifu_bp_hit_taken_q_f) & ~uncacheable_miss_ff ? STREAM : ((((bus_ifu_wr_en_ff & ~exu_flush_final) & ~(bus_ifu_wr_en_ff & last_beat)) & ~ifu_bp_hit_taken_q_f) & ~uncacheable_miss_ff ? STREAM : (((~ic_byp_hit_f & ~exu_flush_final) & (bus_ifu_wr_en_ff & last_beat)) & ~uncacheable_miss_ff ? IDLE : ((exu_flush_final | ifu_bp_hit_taken_q_f) & ~(bus_ifu_wr_en_ff & last_beat) ? HIT_U_MISS : IDLE)))))))));
				miss_state_en = ((((dec_tlu_force_halt | exu_flush_final) | ic_byp_hit_f) | ifu_bp_hit_taken_q_f) | (bus_ifu_wr_en_ff & last_beat)) | (bus_ifu_wr_en_ff & ~uncacheable_miss_ff);
			end
			CRIT_WRD_RDY: begin : crit_wrd_rdy
				miss_nxtstate = IDLE;
				miss_state_en = ((exu_flush_final | flush_final_f) | ic_byp_hit_f) | dec_tlu_force_halt;
			end
			STREAM: begin : stream
				miss_nxtstate = ((((exu_flush_final | ifu_bp_hit_taken_q_f) | stream_eol_f) & ~(bus_ifu_wr_en_ff & last_beat)) & ~dec_tlu_force_halt ? HIT_U_MISS : IDLE);
				miss_state_en = (((exu_flush_final | ifu_bp_hit_taken_q_f) | stream_eol_f) | (bus_ifu_wr_en_ff & last_beat)) | dec_tlu_force_halt;
			end
			MISS_WAIT: begin : miss_wait
				miss_nxtstate = ((exu_flush_final & ~(bus_ifu_wr_en_ff & last_beat)) & ~dec_tlu_force_halt ? HIT_U_MISS : IDLE);
				miss_state_en = (exu_flush_final | (bus_ifu_wr_en_ff & last_beat)) | dec_tlu_force_halt;
			end
			HIT_U_MISS: begin : hit_u_miss
				miss_nxtstate = ((ic_miss_under_miss_f & ~(bus_ifu_wr_en_ff & last_beat)) & ~dec_tlu_force_halt ? SCND_MISS : ((ic_ignore_2nd_miss_f & ~(bus_ifu_wr_en_ff & last_beat)) & ~dec_tlu_force_halt ? STALL_SCND_MISS : IDLE));
				miss_state_en = (((bus_ifu_wr_en_ff & last_beat) | ic_miss_under_miss_f) | ic_ignore_2nd_miss_f) | dec_tlu_force_halt;
			end
			SCND_MISS: begin : scnd_miss
				miss_nxtstate = (dec_tlu_force_halt ? IDLE : (exu_flush_final ? (bus_ifu_wr_en_ff & last_beat ? IDLE : HIT_U_MISS) : CRIT_BYP_OK));
				miss_state_en = ((bus_ifu_wr_en_ff & last_beat) | exu_flush_final) | dec_tlu_force_halt;
			end
			STALL_SCND_MISS: begin : stall_scnd_miss
				miss_nxtstate = (dec_tlu_force_halt ? IDLE : (exu_flush_final ? (bus_ifu_wr_en_ff & last_beat ? IDLE : HIT_U_MISS) : IDLE));
				miss_state_en = ((bus_ifu_wr_en_ff & last_beat) | exu_flush_final) | dec_tlu_force_halt;
			end
			default: begin : def_case
				miss_nxtstate = IDLE;
				miss_state_en = 1'b0;
			end
		endcase
	end
	rvdffs #(.WIDTH(3)) miss_state_ff(
		.clk(active_clk),
		.din(miss_nxtstate),
		.dout({miss_state}),
		.en(miss_state_en),
		.rst_l(rst_l)
	);
	wire sel_hold_imb;
	assign miss_pending = miss_state != IDLE;
	assign crit_wd_byp_ok_ff = (miss_state == CRIT_BYP_OK) | ((miss_state == CRIT_WRD_RDY) & ~flush_final_f);
	assign sel_hold_imb = ((((miss_pending & ~(bus_ifu_wr_en_ff & last_beat)) & ~((miss_state == CRIT_WRD_RDY) & exu_flush_final)) & ~((miss_state == CRIT_WRD_RDY) & crit_byp_hit_f)) | ic_act_miss_f) | (miss_pending & (miss_nxtstate == CRIT_WRD_RDY));
	wire sel_hold_imb_scnd;
	wire [31:1] imb_scnd_in;
	wire [31:1] imb_scnd_ff;
	wire uncacheable_miss_scnd_in;
	wire uncacheable_miss_scnd_ff;
	wire [pt[1060-:7] - 1:0] tagv_mb_scnd_in;
	wire [pt[1060-:7] - 1:0] tagv_mb_scnd_ff;
	wire [pt[1027-:7] - 1:0] way_status_mb_scnd_in;
	wire [pt[1027-:7] - 1:0] way_status_mb_scnd_ff;
	assign sel_hold_imb_scnd = ((miss_state == SCND_MISS) | ic_miss_under_miss_f) & ~flush_final_f;
	assign way_status_mb_scnd_in[pt[1027-:7] - 1:0] = (miss_state == SCND_MISS ? way_status_mb_scnd_ff[pt[1027-:7] - 1:0] : {way_status[pt[1027-:7] - 1:0]});
	assign tagv_mb_scnd_in[pt[1060-:7] - 1:0] = (miss_state == SCND_MISS ? tagv_mb_scnd_ff[pt[1060-:7] - 1:0] : {ic_tag_valid[pt[1060-:7] - 1:0]} & {pt[1060-:7] {~reset_all_tags & ~exu_flush_final}});
	assign uncacheable_miss_scnd_in = (sel_hold_imb_scnd ? uncacheable_miss_scnd_ff : ifc_fetch_uncacheable_bf);
	rvdff_fpga #(.WIDTH(1)) unc_miss_scnd_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din(uncacheable_miss_scnd_in),
		.dout(uncacheable_miss_scnd_ff)
	);
	rvdffpcie #(.WIDTH(31)) imb_f_scnd_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(fetch_bf_f_c1_clken),
		.din({imb_scnd_in[31:1]}),
		.dout({imb_scnd_ff[31:1]})
	);
	rvdff_fpga #(.WIDTH(pt[1027-:7])) mb_rep_wayf2_scnd_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din({way_status_mb_scnd_in[pt[1027-:7] - 1:0]}),
		.dout({way_status_mb_scnd_ff[pt[1027-:7] - 1:0]})
	);
	rvdff_fpga #(.WIDTH(pt[1060-:7])) mb_tagv_scnd_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din({tagv_mb_scnd_in[pt[1060-:7] - 1:0]}),
		.dout({tagv_mb_scnd_ff[pt[1060-:7] - 1:0]})
	);
	assign ic_req_addr_bits_hi_3[pt[1182-:8]:3] = bus_rd_addr_count[pt[1174-:8] - 1:0];
	assign ic_wr_addr_bits_hi_3[pt[1182-:8]:3] = ifu_bus_rid_ff[pt[1174-:8] - 1:0] & {pt[1174-:8] {bus_ifu_wr_en_ff}};
	assign fetch_req_icache_f = (ifc_fetch_req_f & ~ifc_iccm_access_f) & ~ifc_region_acc_fault_final_f;
	assign fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f;
	assign ic_iccm_hit_f = fetch_req_iccm_f & ((~miss_pending | (miss_state == HIT_U_MISS)) | (miss_state == STREAM));
	assign ic_byp_hit_f = ((crit_byp_hit_f | stream_hit_f) & fetch_req_icache_f) & miss_pending;
	assign ic_act_hit_f = (((|ic_rd_hit[pt[1060-:7] - 1:0] & fetch_req_icache_f) & ~reset_all_tags) & (~miss_pending | (miss_state == HIT_U_MISS))) & ~sel_mb_addr_ff;
	assign ic_act_miss_f = ((((~(|ic_rd_hit[pt[1060-:7] - 1:0]) | reset_all_tags) & fetch_req_icache_f) & ~miss_pending) | scnd_miss_req) & ~ifc_region_acc_fault_final_f;
	assign ic_miss_under_miss_f = ((((((~(|ic_rd_hit[pt[1060-:7] - 1:0]) | reset_all_tags) & fetch_req_icache_f) & (miss_state == HIT_U_MISS)) & (imb_ff[31:pt[998-:7]] != ifu_fetch_addr_int_f[31:pt[998-:7]])) & ~uncacheable_miss_ff) & ~sel_mb_addr_ff) & ~ifc_region_acc_fault_final_f;
	assign ic_ignore_2nd_miss_f = (((~(|ic_rd_hit[pt[1060-:7] - 1:0]) | reset_all_tags) & fetch_req_icache_f) & (miss_state == HIT_U_MISS)) & ((imb_ff[31:pt[998-:7]] == ifu_fetch_addr_int_f[31:pt[998-:7]]) | uncacheable_miss_ff);
	assign ic_hit_f = ((ic_act_hit_f | ic_byp_hit_f) | ic_iccm_hit_f) | (ifc_region_acc_fault_final_f & ifc_fetch_req_f);
	assign uncacheable_miss_in = (scnd_miss_req ? uncacheable_miss_scnd_ff : (sel_hold_imb ? uncacheable_miss_ff : ifc_fetch_uncacheable_bf));
	assign imb_in[31:1] = (scnd_miss_req ? imb_scnd_ff[31:1] : (sel_hold_imb ? imb_ff[31:1] : {ifc_fetch_addr_bf[31:1]}));
	assign imb_scnd_in[31:1] = (sel_hold_imb_scnd ? imb_scnd_ff[31:1] : {ifc_fetch_addr_bf[31:1]});
	assign scnd_miss_index_match = ((imb_ff[pt[1104-:9]:pt[998-:7]] == imb_scnd_ff[pt[1104-:9]:pt[998-:7]]) & scnd_miss_req) & ~ifu_wr_cumulative_err_data;
	assign way_status_mb_in[pt[1027-:7] - 1:0] = (scnd_miss_req & ~scnd_miss_index_match ? way_status_mb_scnd_ff[pt[1027-:7] - 1:0] : (scnd_miss_req & scnd_miss_index_match ? way_status_rep_new[pt[1027-:7] - 1:0] : (miss_pending ? way_status_mb_ff[pt[1027-:7] - 1:0] : {way_status[pt[1027-:7] - 1:0]})));
	assign tagv_mb_in[pt[1060-:7] - 1:0] = (scnd_miss_req ? tagv_mb_scnd_ff[pt[1060-:7] - 1:0] | ({pt[1060-:7] {scnd_miss_index_match}} & replace_way_mb_any[pt[1060-:7] - 1:0]) : (miss_pending ? tagv_mb_ff[pt[1060-:7] - 1:0] : {ic_tag_valid[pt[1060-:7] - 1:0]} & {pt[1060-:7] {~reset_all_tags & ~exu_flush_final}}));
	assign reset_ic_in = (miss_pending & ~scnd_miss_req_q) & (reset_all_tags | reset_ic_ff);
	rvdffpcie #(.WIDTH(31)) ifu_fetch_addr_f_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(fetch_bf_f_c1_clken),
		.din({ifc_fetch_addr_bf[31:1]}),
		.dout({ifu_fetch_addr_int_f[31:1]})
	);
	assign vaddr_f[pt[1182-:8]:1] = ifu_fetch_addr_int_f[pt[1182-:8]:1];
	rvdffpcie #(.WIDTH(31)) imb_f_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(fetch_bf_f_c1_clken),
		.din(imb_in[31:1]),
		.dout(imb_ff[31:1])
	);
	rvdff_fpga #(.WIDTH(1)) unc_miss_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din(uncacheable_miss_in),
		.dout(uncacheable_miss_ff)
	);
	assign miss_addr_in[31:pt[1182-:8] + 1] = (~miss_pending ? imb_ff[31:pt[1182-:8] + 1] : (scnd_miss_req_q ? imb_scnd_ff[31:pt[1182-:8] + 1] : miss_addr[31:pt[1182-:8] + 1]));
	rvdfflie #(
		.WIDTH(31 - pt[1182-:8]),
		.LEFT((31 - pt[1182-:8]) - 8)
	) miss_f_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en((bus_ifu_bus_clk_en | ic_act_miss_f) | dec_tlu_force_halt),
		.din({miss_addr_in[31:pt[1182-:8] + 1]}),
		.dout({miss_addr[31:pt[1182-:8] + 1]})
	);
	rvdff_fpga #(.WIDTH(pt[1027-:7])) mb_rep_wayf2_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din({way_status_mb_in[pt[1027-:7] - 1:0]}),
		.dout({way_status_mb_ff[pt[1027-:7] - 1:0]})
	);
	rvdff_fpga #(.WIDTH(pt[1060-:7])) mb_tagv_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din({tagv_mb_in[pt[1060-:7] - 1:0]}),
		.dout({tagv_mb_ff[pt[1060-:7] - 1:0]})
	);
	assign ifc_fetch_req_qual_bf = (ifc_fetch_req_bf & ~((miss_state == CRIT_WRD_RDY) & flush_final_f)) & ~stream_miss_f;
	assign ifc_fetch_req_f = ifc_fetch_req_f_raw & ~exu_flush_final;
	rvdff_fpga #(.WIDTH(1)) ifu_iccm_acc_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din(ifc_iccm_access_bf),
		.dout(ifc_iccm_access_f)
	);
	rvdff_fpga #(.WIDTH(1)) ifu_iccm_reg_acc_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din(ifc_region_acc_fault_final_bf),
		.dout(ifc_region_acc_fault_final_f)
	);
	rvdff_fpga #(.WIDTH(1)) rgn_acc_ff(
		.rst_l(rst_l),
		.clk(fetch_bf_f_c1_clk),
		.clken(fetch_bf_f_c1_clken),
		.rawclk(clk),
		.din(ifc_region_acc_fault_bf),
		.dout(ifc_region_acc_fault_f)
	);
	assign ifu_ic_req_addr_f[31:3] = {miss_addr[31:pt[1182-:8] + 1], ic_req_addr_bits_hi_3[pt[1182-:8]:3]};
	assign ifu_ic_mb_empty = (((miss_state == HIT_U_MISS) | (miss_state == STREAM)) & ~(bus_ifu_wr_en_ff & last_beat)) | ~miss_pending;
	assign ifu_miss_state_idle = miss_state == IDLE;
	assign sel_mb_addr = ((miss_pending & write_ic_16_bytes) & ~uncacheable_miss_ff) | reset_tag_valid_for_miss;
	assign ifu_ic_rw_int_addr[31:1] = ({31 {sel_mb_addr}} & {imb_ff[31:pt[1182-:8] + 1], ic_wr_addr_bits_hi_3[pt[1182-:8]:3], imb_ff[2:1]}) | ({31 {~sel_mb_addr}} & ifc_fetch_addr_bf[31:1]);
	assign sel_mb_status_addr = ((((miss_pending & write_ic_16_bytes) & ~uncacheable_miss_ff) & last_beat) & bus_ifu_wr_en_ff_q) | reset_tag_valid_for_miss;
	assign ifu_status_wr_addr[31:1] = ({31 {sel_mb_status_addr}} & {imb_ff[31:pt[1182-:8] + 1], ic_wr_addr_bits_hi_3[pt[1182-:8]:3], imb_ff[2:1]}) | ({31 {~sel_mb_status_addr}} & ifu_fetch_addr_int_f[31:1]);
	assign ic_rw_addr[31:1] = ifu_ic_rw_int_addr[31:1];
	generate
		if (pt[1125-:5] == 1) begin : icache_ecc_1
			wire [6:0] ic_wr_ecc;
			wire [6:0] ic_miss_buff_ecc;
			wire [141:0] ic_wr_16bytes_data;
			wire [70:0] ifu_ic_debug_rd_data_in;
			rvecc_encode_64 ic_ecc_encode_64_bus(
				.din(ifu_bus_rdata_ff[63:0]),
				.ecc_out(ic_wr_ecc[6:0])
			);
			rvecc_encode_64 ic_ecc_encode_64_buff(
				.din(ic_miss_buff_half[63:0]),
				.ecc_out(ic_miss_buff_ecc[6:0])
			);
			genvar i;
			for (i = 0; i < pt[1189-:7]; i = i + 1) begin : ic_wr_data_loop
				assign ic_wr_data[(i * 71) + 70-:71] = ic_wr_16bytes_data[(71 * i) + 70:71 * i];
			end
			assign ic_debug_wr_data[70:0] = {dec_tlu_ic_diag_pkt[89:19]};
			assign ic_error_start = (|ic_eccerr[pt[1189-:7] - 1:0] & ic_act_hit_f) | ic_rd_parity_final_err;
			assign ifu_ic_debug_rd_data_in[70:0] = (ic_debug_ict_array_sel_ff ? {2'b00, ictag_debug_rd_data[25:21], 32'b00000000000000000000000000000000, ictag_debug_rd_data[20:0], {7 - pt[1027-:7] {1'b0}}, way_status[pt[1027-:7] - 1:0], 3'b000, ic_debug_tag_val_rd_out} : ic_debug_rd_data[70:0]);
			rvdffe #(.WIDTH(71)) ifu_debug_data_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(debug_data_clken),
				.din({ifu_ic_debug_rd_data_in[70:0]}),
				.dout({ifu_ic_debug_rd_data[70:0]})
			);
			assign ic_wr_16bytes_data[141:0] = (ifu_bus_rid_ff[0] ? {ic_wr_ecc[6:0], ifu_bus_rdata_ff[63:0], ic_miss_buff_ecc[6:0], ic_miss_buff_half[63:0]} : {ic_miss_buff_ecc[6:0], ic_miss_buff_half[63:0], ic_wr_ecc[6:0], ifu_bus_rdata_ff[63:0]});
		end
		else begin : icache_parity_1
			wire [3:0] ic_wr_parity;
			wire [3:0] ic_miss_buff_parity;
			wire [135:0] ic_wr_16bytes_data;
			wire [70:0] ifu_ic_debug_rd_data_in;
			genvar i;
			for (i = 0; i < 4; i = i + 1) begin : DATA_PGEN
				rveven_paritygen #(.WIDTH(16)) par_bus(
					.data_in(ifu_bus_rdata_ff[(16 * i) + 15:16 * i]),
					.parity_out(ic_wr_parity[i])
				);
				rveven_paritygen #(.WIDTH(16)) par_buff(
					.data_in(ic_miss_buff_half[(16 * i) + 15:16 * i]),
					.parity_out(ic_miss_buff_parity[i])
				);
			end
			for (i = 0; i < pt[1189-:7]; i = i + 1) begin : ic_wr_data_loop
				assign ic_wr_data[(i * 71) + 70-:71] = {3'b000, ic_wr_16bytes_data[(68 * i) + 67:68 * i]};
			end
			assign ic_debug_wr_data[70:0] = {dec_tlu_ic_diag_pkt[89:19]};
			assign ic_error_start = (|ic_parerr[pt[1189-:7] - 1:0] & ic_act_hit_f) | ic_rd_parity_final_err;
			assign ifu_ic_debug_rd_data_in[70:0] = (ic_debug_ict_array_sel_ff ? {6'b000000, ictag_debug_rd_data[21], 32'b00000000000000000000000000000000, ictag_debug_rd_data[20:0], {7 - pt[1027-:7] {1'b0}}, way_status[pt[1027-:7] - 1:0], 3'b000, ic_debug_tag_val_rd_out} : ic_debug_rd_data[70:0]);
			rvdffe #(.WIDTH(71)) ifu_debug_data_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(debug_data_clken),
				.din({ifu_ic_debug_rd_data_in[70:0]}),
				.dout({ifu_ic_debug_rd_data[70:0]})
			);
			assign ic_wr_16bytes_data[135:0] = (ifu_bus_rid_ff[0] ? {ic_wr_parity[3:0], ifu_bus_rdata_ff[63:0], ic_miss_buff_parity[3:0], ic_miss_buff_half[63:0]} : {ic_miss_buff_parity[3:0], ic_miss_buff_half[63:0], ic_wr_parity[3:0], ifu_bus_rdata_ff[63:0]});
		end
	endgenerate
	assign ifu_wr_data_comb_err = bus_ifu_wr_data_error_ff;
	assign ifu_wr_cumulative_err = (ifu_wr_data_comb_err | ifu_wr_data_comb_err_ff) & ~reset_beat_cnt;
	assign ifu_wr_cumulative_err_data = ifu_wr_data_comb_err | ifu_wr_data_comb_err_ff;
	assign sel_byp_data = (ic_crit_wd_rdy | (miss_state == STREAM)) | (miss_state == CRIT_BYP_OK);
	assign sel_ic_data = (~(((ic_crit_wd_rdy | (miss_state == STREAM)) | (miss_state == CRIT_BYP_OK)) | (miss_state == MISS_WAIT)) & ~fetch_req_iccm_f) & ~ifc_region_acc_fault_final_f;
	generate
		if (pt[922-:5] == 1) begin : iccm_icache
			assign sel_iccm_data = fetch_req_iccm_f;
			assign ic_final_data[63:0] = {64 {(sel_byp_data | sel_iccm_data) | sel_ic_data}} & {ic_rd_data[63:0]};
			assign ic_premux_data[63:0] = ({64 {sel_byp_data}} & {ic_byp_data_only_new[63:0]}) | ({64 {sel_iccm_data}} & {iccm_rd_data[63:0]});
			assign ic_sel_premux_data = sel_iccm_data | sel_byp_data;
		end
	endgenerate
	generate
		if (pt[900-:5] == 1) begin : iccm_only
			assign sel_iccm_data = fetch_req_iccm_f;
			assign ic_final_data[63:0] = ({64 {sel_byp_data}} & {ic_byp_data_only_new[63:0]}) | ({64 {sel_iccm_data}} & {iccm_rd_data[63:0]});
			assign ic_premux_data = {64 {1'sb0}};
			assign ic_sel_premux_data = 1'b0;
		end
	endgenerate
	generate
		if (pt[1053-:5] == 1) begin : icache_only
			assign ic_final_data[63:0] = {64 {sel_byp_data | sel_ic_data}} & {ic_rd_data[63:0]};
			assign ic_premux_data[63:0] = {64 {sel_byp_data}} & {ic_byp_data_only_new[63:0]};
			assign ic_sel_premux_data = sel_byp_data;
		end
	endgenerate
	generate
		if (pt[140-:5] == 1) begin : no_iccm_no_icache
			assign ic_final_data[63:0] = {64 {sel_byp_data}} & {ic_byp_data_only_new[63:0]};
			assign ic_premux_data = 0;
			assign ic_sel_premux_data = 1'b0;
		end
	endgenerate
	assign ifc_bus_acc_fault_f[1:0] = {2 {ic_byp_hit_f}} & ifu_byp_data_err_f[1:0];
	assign ic_data_f[31:0] = ic_final_data[31:0];
	assign fetch_req_f_qual = ic_hit_f & ~exu_flush_final;
	assign ic_access_fault_f[1:0] = ({2 {ifc_region_acc_fault_final_f}} | ifc_bus_acc_fault_f[1:0]) & {2 {~exu_flush_final}};
	assign ic_access_fault_type_f[1:0] = (|iccm_rd_ecc_double_err ? 2'b01 : (ifc_region_acc_fault_f ? 2'b10 : (ifc_region_acc_fault_memory_f ? 2'b11 : 2'b00)));
	localparam [1:0] ERR_FETCH2 = 2'b10;
	assign ic_fetch_val_f[1] = ((fetch_req_f_qual & ifu_bp_inst_mask_f) & ~(vaddr_f[pt[1182-:8]:1] == {pt[1182-:8] {1'b1}})) & (err_stop_state != ERR_FETCH2);
	assign ic_fetch_val_f[0] = fetch_req_f_qual;
	assign two_byte_instr = ic_data_f[1:0] != 2'b11;
	wire [63:0] ic_miss_buff_data_in;
	assign ic_miss_buff_data_in[63:0] = ifu_bus_rsp_rdata[63:0];
	generate
		genvar i;
		for (i = 0; i < pt[1084-:8]; i = i + 1) begin : wr_flop
			function automatic signed [pt[826-:8] - 1:0] sv2v_cast_ADFF4_signed;
				input reg signed [pt[826-:8] - 1:0] inp;
				sv2v_cast_ADFF4_signed = inp;
			endfunction
			assign write_fill_data[i] = bus_ifu_wr_en & (sv2v_cast_ADFF4_signed(i) == ifu_bus_rsp_tag[pt[826-:8] - 1:0]);
			rvdffe #(.WIDTH(32)) byp_data_0_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(write_fill_data[i]),
				.din(ic_miss_buff_data_in[31:0]),
				.dout(ic_miss_buff_data[((i * 2) * 32) + 31-:32])
			);
			rvdffe #(.WIDTH(32)) byp_data_1_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.en(write_fill_data[i]),
				.din(ic_miss_buff_data_in[63:32]),
				.dout(ic_miss_buff_data[(((i * 2) + 1) * 32) + 31-:32])
			);
			assign ic_miss_buff_data_valid_in[i] = (write_fill_data[i] ? 1'b1 : ic_miss_buff_data_valid[i] & ~ic_act_miss_f);
			rvdff #(.WIDTH(1)) byp_data_valid_ff(
				.rst_l(rst_l),
				.clk(active_clk),
				.din(ic_miss_buff_data_valid_in[i]),
				.dout(ic_miss_buff_data_valid[i])
			);
			assign ic_miss_buff_data_error_in[i] = (write_fill_data[i] ? bus_ifu_wr_data_error : ic_miss_buff_data_error[i] & ~ic_act_miss_f);
			rvdff #(.WIDTH(1)) byp_data_error_ff(
				.rst_l(rst_l),
				.clk(active_clk),
				.din(ic_miss_buff_data_error_in[i]),
				.dout(ic_miss_buff_data_error[i])
			);
		end
	endgenerate
	wire [pt[1182-:8]:1] bypass_index;
	wire [pt[1182-:8]:3] bypass_index_5_3_inc;
	wire bypass_data_ready_in;
	wire ic_crit_wd_rdy_new_in;
	assign bypass_index[pt[1182-:8]:1] = imb_ff[pt[1182-:8]:1];
	assign bypass_index_5_3_inc[pt[1182-:8]:3] = bypass_index[pt[1182-:8]:3] + 1;
	assign bypass_data_ready_in = (((((ic_miss_buff_data_valid_in[bypass_index[pt[1182-:8]:3]] & ~bypass_index[2]) & ~bypass_index[1]) | ((ic_miss_buff_data_valid_in[bypass_index[pt[1182-:8]:3]] & ~bypass_index[2]) & bypass_index[1])) | ((ic_miss_buff_data_valid_in[bypass_index[pt[1182-:8]:3]] & bypass_index[2]) & ~bypass_index[1])) | (((ic_miss_buff_data_valid_in[bypass_index[pt[1182-:8]:3]] & ic_miss_buff_data_valid_in[bypass_index_5_3_inc[pt[1182-:8]:3]]) & bypass_index[2]) & bypass_index[1])) | (ic_miss_buff_data_valid_in[bypass_index[pt[1182-:8]:3]] & (bypass_index[pt[1182-:8]:3] == {pt[1182-:8] {1'b1}}));
	assign ic_crit_wd_rdy_new_in = (((((bypass_data_ready_in & crit_wd_byp_ok_ff) & uncacheable_miss_ff) & ~exu_flush_final) & ~ifu_bp_hit_taken_q_f) | (((crit_wd_byp_ok_ff & ~uncacheable_miss_ff) & ~exu_flush_final) & ~ifu_bp_hit_taken_q_f)) | (((ic_crit_wd_rdy_new_ff & ~fetch_req_icache_f) & crit_wd_byp_ok_ff) & ~exu_flush_final);
	assign byp_fetch_index[pt[1182-:8]:1] = ifu_fetch_addr_int_f[pt[1182-:8]:1];
	assign byp_fetch_index_0[pt[1182-:8]:2] = {ifu_fetch_addr_int_f[pt[1182-:8]:3], 1'b0};
	assign byp_fetch_index_1[pt[1182-:8]:2] = {ifu_fetch_addr_int_f[pt[1182-:8]:3], 1'b1};
	assign byp_fetch_index_inc[pt[1182-:8]:3] = ifu_fetch_addr_int_f[pt[1182-:8]:3] + 1'b1;
	assign byp_fetch_index_inc_0[pt[1182-:8]:2] = {byp_fetch_index_inc[pt[1182-:8]:3], 1'b0};
	assign byp_fetch_index_inc_1[pt[1182-:8]:2] = {byp_fetch_index_inc[pt[1182-:8]:3], 1'b1};
	assign ifu_byp_data_err_new = ((((~ifu_fetch_addr_int_f[2] & ~ifu_fetch_addr_int_f[1]) & ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]]) | ((~ifu_fetch_addr_int_f[2] & ifu_fetch_addr_int_f[1]) & ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]])) | ((ifu_fetch_addr_int_f[2] & ~ifu_fetch_addr_int_f[1]) & ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]])) | ((ifu_fetch_addr_int_f[2] & ifu_fetch_addr_int_f[1]) & (ic_miss_buff_data_error[byp_fetch_index_inc[pt[1182-:8]:3]] | ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]]));
	assign ifu_byp_data_err_f[1:0] = (ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]] ? 2'b11 : (((ifu_fetch_addr_int_f[2] & ifu_fetch_addr_int_f[1]) & ~ic_miss_buff_data_error[byp_fetch_index[pt[1182-:8]:3]]) & (~miss_wrap_f & ic_miss_buff_data_error[byp_fetch_index_inc[pt[1182-:8]:3]]) ? 2'b10 : 2'b00));
	assign ic_byp_data_only_pre_new[79:0] = ({80 {~ifu_fetch_addr_int_f[2]}} & {ic_miss_buff_data[(byp_fetch_index_inc_0 * 32) + 15-:16], ic_miss_buff_data[(byp_fetch_index_1 * 32) + 31-:32], ic_miss_buff_data[(byp_fetch_index_0 * 32) + 31-:32]}) | ({80 {ifu_fetch_addr_int_f[2]}} & {ic_miss_buff_data[(byp_fetch_index_inc_1 * 32) + 15-:16], ic_miss_buff_data[(byp_fetch_index_inc_0 * 32) + 31-:32], ic_miss_buff_data[(byp_fetch_index_1 * 32) + 31-:32]});
	assign ic_byp_data_only_new[79:0] = (~ifu_fetch_addr_int_f[1] ? {ic_byp_data_only_pre_new[79:0]} : {16'b0000000000000000, ic_byp_data_only_pre_new[79:16]});
	assign miss_wrap_f = imb_ff[pt[998-:7]] != ifu_fetch_addr_int_f[pt[998-:7]];
	assign miss_buff_hit_unq_f = (((((ic_miss_buff_data_valid[byp_fetch_index[pt[1182-:8]:3]] & ~byp_fetch_index[2]) & ~byp_fetch_index[1]) | ((ic_miss_buff_data_valid[byp_fetch_index[pt[1182-:8]:3]] & ~byp_fetch_index[2]) & byp_fetch_index[1])) | ((ic_miss_buff_data_valid[byp_fetch_index[pt[1182-:8]:3]] & byp_fetch_index[2]) & ~byp_fetch_index[1])) | (((ic_miss_buff_data_valid[byp_fetch_index[pt[1182-:8]:3]] & ic_miss_buff_data_valid[byp_fetch_index_inc[pt[1182-:8]:3]]) & byp_fetch_index[2]) & byp_fetch_index[1])) | (ic_miss_buff_data_valid[byp_fetch_index[pt[1182-:8]:3]] & (byp_fetch_index[pt[1182-:8]:3] == {pt[1174-:8] {1'b1}}));
	assign stream_hit_f = (miss_buff_hit_unq_f & ~miss_wrap_f) & (miss_state == STREAM);
	assign stream_miss_f = (~(miss_buff_hit_unq_f & ~miss_wrap_f) & (miss_state == STREAM)) & ifc_fetch_req_f;
	assign stream_eol_f = ((byp_fetch_index[pt[1182-:8]:2] == {pt[1174-:8] + 1 {1'b1}}) & ifc_fetch_req_f) & stream_hit_f;
	assign crit_byp_hit_f = miss_buff_hit_unq_f & ((miss_state == CRIT_WRD_RDY) | (miss_state == CRIT_BYP_OK));
	assign other_tag[pt[826-:8] - 1:0] = {ifu_bus_rid_ff[pt[826-:8] - 1:1], ~ifu_bus_rid_ff[0]};
	assign second_half_available = ic_miss_buff_data_valid[other_tag];
	assign write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff;
	assign ic_miss_buff_half[63:0] = {ic_miss_buff_data[{other_tag, 1'b1} * 32+:32], ic_miss_buff_data[{other_tag, 1'b0} * 32+:32]};
	assign ic_rd_parity_final_err = (((ic_tag_perr & ~exu_flush_final) & sel_ic_data) & ~(ifc_region_acc_fault_final_f | |ifc_bus_acc_fault_f)) & (((fetch_req_icache_f & ~reset_all_tags) & (~miss_pending | (miss_state == HIT_U_MISS))) & ~sel_mb_addr_ff);
	wire [pt[1060-:7] - 1:0] perr_err_inv_way;
	wire [pt[1104-:9]:pt[998-:7]] perr_ic_index_ff;
	reg perr_sel_invalidate;
	reg perr_sb_write_status;
	rvdffe #(
		.WIDTH((pt[1104-:9] - pt[998-:7]) + 1),
		.OVERRIDE(1)
	) perr_dat_ff(
		.din(ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7]]),
		.dout(perr_ic_index_ff[pt[1104-:9]:pt[998-:7]]),
		.en(perr_sb_write_status),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	assign perr_err_inv_way[pt[1060-:7] - 1:0] = {pt[1060-:7] {perr_sel_invalidate}};
	localparam [2:0] ECC_CORR = 3'b011;
	assign iccm_correct_ecc = perr_state == ECC_CORR;
	assign dma_sb_err_state = perr_state == DMA_SB_ERR;
	assign iccm_buf_correct_ecc = iccm_correct_ecc & ~dma_sb_err_state_ff;
	localparam [2:0] ECC_WFF = 3'b010;
	localparam [2:0] ERR_IDLE = 3'b000;
	localparam [2:0] IC_WFF = 3'b001;
	always @(*) begin : ERROR_SM
		perr_nxtstate = ERR_IDLE;
		perr_state_en = 1'b0;
		perr_sb_write_status = 1'b0;
		perr_sel_invalidate = 1'b0;
		case (perr_state)
			ERR_IDLE: begin : err_idle
				perr_nxtstate = (iccm_dma_sb_error ? DMA_SB_ERR : (ic_error_start & ~exu_flush_final ? IC_WFF : ECC_WFF));
				perr_state_en = (((iccm_error_start | ic_error_start) & ~exu_flush_final) | iccm_dma_sb_error) & ~dec_tlu_force_halt;
				perr_sb_write_status = perr_state_en;
			end
			IC_WFF: begin : icache_wff
				perr_nxtstate = ERR_IDLE;
				perr_state_en = dec_tlu_flush_lower_wb | dec_tlu_force_halt;
				perr_sel_invalidate = dec_tlu_flush_err_wb & dec_tlu_flush_lower_wb;
			end
			ECC_WFF: begin : ecc_wff
				perr_nxtstate = ((~dec_tlu_flush_err_wb & dec_tlu_flush_lower_wb) | dec_tlu_force_halt ? ERR_IDLE : ECC_CORR);
				perr_state_en = dec_tlu_flush_lower_wb | dec_tlu_force_halt;
			end
			DMA_SB_ERR: begin : dma_sb_ecc
				perr_nxtstate = (dec_tlu_force_halt ? ERR_IDLE : ECC_CORR);
				perr_state_en = 1'b1;
			end
			ECC_CORR: begin : ecc_corr
				perr_nxtstate = ERR_IDLE;
				perr_state_en = 1'b1;
			end
			default: begin : def_case
				perr_nxtstate = ERR_IDLE;
				perr_state_en = 1'b0;
				perr_sb_write_status = 1'b0;
				perr_sel_invalidate = 1'b0;
			end
		endcase
	end
	rvdffs #(.WIDTH(3)) perr_state_ff(
		.clk(active_clk),
		.din(perr_nxtstate),
		.dout({perr_state}),
		.en(perr_state_en),
		.rst_l(rst_l)
	);
	localparam [1:0] ERR_FETCH1 = 2'b01;
	localparam [1:0] ERR_STOP_IDLE = 2'b00;
	always @(*) begin : ERROR_STOP_FETCH
		err_stop_nxtstate = ERR_STOP_IDLE;
		err_stop_state_en = 1'b0;
		err_stop_fetch = 1'b0;
		iccm_correction_state = 1'b0;
		case (err_stop_state)
			ERR_STOP_IDLE: begin : err_stop_idle
				err_stop_nxtstate = ERR_FETCH1;
				err_stop_state_en = (dec_tlu_flush_err_wb & (perr_state == ECC_WFF)) & ~dec_tlu_force_halt;
			end
			ERR_FETCH1: begin : err_fetch1
				err_stop_nxtstate = ((dec_tlu_flush_lower_wb | dec_tlu_i0_commit_cmt) | dec_tlu_force_halt ? ERR_STOP_IDLE : ((ifu_fetch_val[1:0] == 2'b11) | (ifu_fetch_val[0] & two_byte_instr) ? ERR_STOP_FETCH : (ifu_fetch_val[0] ? ERR_FETCH2 : ERR_FETCH1)));
				err_stop_state_en = (((dec_tlu_flush_lower_wb | dec_tlu_i0_commit_cmt) | ifu_fetch_val[0]) | ifu_bp_hit_taken_q_f) | dec_tlu_force_halt;
				err_stop_fetch = ((ifu_fetch_val[1:0] == 2'b11) | (ifu_fetch_val[0] & two_byte_instr)) & ~(exu_flush_final | dec_tlu_i0_commit_cmt);
				iccm_correction_state = 1'b1;
			end
			ERR_FETCH2: begin : err_fetch2
				err_stop_nxtstate = ((dec_tlu_flush_lower_wb | dec_tlu_i0_commit_cmt) | dec_tlu_force_halt ? ERR_STOP_IDLE : (ifu_fetch_val[0] ? ERR_STOP_FETCH : ERR_FETCH2));
				err_stop_state_en = ((dec_tlu_flush_lower_wb | dec_tlu_i0_commit_cmt) | ifu_fetch_val[0]) | dec_tlu_force_halt;
				err_stop_fetch = (ifu_fetch_val[0] & ~exu_flush_final) & ~dec_tlu_i0_commit_cmt;
				iccm_correction_state = 1'b1;
			end
			ERR_STOP_FETCH: begin : ecc_wff
				err_stop_nxtstate = (((dec_tlu_flush_lower_wb & ~dec_tlu_flush_err_wb) | dec_tlu_i0_commit_cmt) | dec_tlu_force_halt ? ERR_STOP_IDLE : (dec_tlu_flush_err_wb ? ERR_FETCH1 : ERR_STOP_FETCH));
				err_stop_state_en = (dec_tlu_flush_lower_wb | dec_tlu_i0_commit_cmt) | dec_tlu_force_halt;
				err_stop_fetch = 1'b1;
				iccm_correction_state = 1'b1;
			end
			default: begin : def_case
				err_stop_nxtstate = ERR_STOP_IDLE;
				err_stop_state_en = 1'b0;
				err_stop_fetch = 1'b0;
				iccm_correction_state = 1'b1;
			end
		endcase
	end
	rvdffs #(.WIDTH(2)) err_stop_state_ff(
		.clk(active_clk),
		.din(err_stop_nxtstate),
		.dout({err_stop_state}),
		.en(err_stop_state_en),
		.rst_l(rst_l)
	);
	assign bus_ifu_bus_clk_en = ifu_bus_clk_en;
	rvclkhdr bus_clk_f(
		.en(bus_ifu_bus_clk_en),
		.l1clk(busclk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr bus_clk(
		.en(bus_ifu_bus_clk_en | dec_tlu_force_halt),
		.l1clk(busclk_force),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign scnd_miss_req = scnd_miss_req_q & ~exu_flush_final;
	assign ifc_bus_ic_req_ff_in = (((ic_act_miss_f | bus_cmd_req_hold) | ifu_bus_cmd_valid) & ~dec_tlu_force_halt) & ~((((bus_cmd_beat_count == {pt[1174-:8] {1'b1}}) & ifu_bus_cmd_valid) & ifu_bus_cmd_ready) & miss_pending);
	rvdff_fpga #(.WIDTH(1)) bus_ic_req_ff2(
		.rst_l(rst_l),
		.clk(busclk_force),
		.clken(bus_ifu_bus_clk_en | dec_tlu_force_halt),
		.rawclk(clk),
		.din(ifc_bus_ic_req_ff_in),
		.dout(ifu_bus_cmd_valid)
	);
	assign bus_cmd_req_in = ((ic_act_miss_f | bus_cmd_req_hold) & ~bus_cmd_sent) & ~dec_tlu_force_halt;
	assign ifu_axi_arvalid = ifu_bus_cmd_valid;
	function automatic [pt[826-:8] - 1:0] sv2v_cast_ADFF4;
		input reg [pt[826-:8] - 1:0] inp;
		sv2v_cast_ADFF4 = inp;
	endfunction
	assign ifu_axi_arid[pt[826-:8] - 1:0] = sv2v_cast_ADFF4(bus_rd_addr_count[pt[1174-:8] - 1:0]) & {pt[826-:8] {ifu_bus_cmd_valid}};
	assign ifu_axi_araddr[31:0] = {ifu_ic_req_addr_f[31:3], 3'b000} & {32 {ifu_bus_cmd_valid}};
	assign ifu_axi_arsize[2:0] = 3'b011;
	assign ifu_axi_arprot[2:0] = 3'b101;
	assign ifu_axi_arcache[3:0] = 4'b1111;
	assign ifu_axi_arregion[3:0] = ifu_ic_req_addr_f[31:28];
	assign ifu_axi_arlen[7:0] = {8 {1'sb0}};
	assign ifu_axi_arburst[1:0] = 2'b01;
	assign ifu_axi_arqos[3:0] = {4 {1'sb0}};
	assign ifu_axi_arlock = 1'b0;
	assign ifu_axi_rready = 1'b1;
	assign ifu_axi_awvalid = 1'b0;
	assign ifu_axi_awid[pt[826-:8] - 1:0] = {pt[826-:8] {1'sb0}};
	assign ifu_axi_awaddr[31:0] = {32 {1'sb0}};
	assign ifu_axi_awsize[2:0] = {3 {1'sb0}};
	assign ifu_axi_awprot[2:0] = {3 {1'sb0}};
	assign ifu_axi_awcache[3:0] = {4 {1'sb0}};
	assign ifu_axi_awregion[3:0] = {4 {1'sb0}};
	assign ifu_axi_awlen[7:0] = {8 {1'sb0}};
	assign ifu_axi_awburst[1:0] = {2 {1'sb0}};
	assign ifu_axi_awqos[3:0] = {4 {1'sb0}};
	assign ifu_axi_awlock = 1'b0;
	assign ifu_axi_wvalid = 1'b0;
	assign ifu_axi_wstrb[7:0] = {8 {1'sb0}};
	assign ifu_axi_wdata[63:0] = {64 {1'sb0}};
	assign ifu_axi_wlast = 1'b0;
	assign ifu_axi_bready = 1'b0;
	assign ifu_bus_arready_unq = ifu_axi_arready;
	assign ifu_bus_rvalid_unq = ifu_axi_rvalid;
	assign ifu_bus_arvalid = ifu_axi_arvalid;
	rvdff_fpga #(.WIDTH(1)) bus_rdy_ff(
		.rst_l(rst_l),
		.clk(busclk),
		.clken(bus_ifu_bus_clk_en),
		.rawclk(clk),
		.din(ifu_bus_arready_unq),
		.dout(ifu_bus_arready_unq_ff)
	);
	rvdff_fpga #(.WIDTH(1)) bus_rsp_vld_ff(
		.rst_l(rst_l),
		.clk(busclk),
		.clken(bus_ifu_bus_clk_en),
		.rawclk(clk),
		.din(ifu_bus_rvalid_unq),
		.dout(ifu_bus_rvalid_unq_ff)
	);
	rvdff_fpga #(.WIDTH(1)) bus_cmd_ff(
		.rst_l(rst_l),
		.clk(busclk),
		.clken(bus_ifu_bus_clk_en),
		.rawclk(clk),
		.din(ifu_bus_arvalid),
		.dout(ifu_bus_arvalid_ff)
	);
	rvdff_fpga #(.WIDTH(2)) bus_rsp_cmd_ff(
		.rst_l(rst_l),
		.clk(busclk),
		.clken(bus_ifu_bus_clk_en),
		.rawclk(clk),
		.din(ifu_axi_rresp[1:0]),
		.dout(ifu_bus_rresp_ff[1:0])
	);
	rvdff_fpga #(.WIDTH(pt[826-:8])) bus_rsp_tag_ff(
		.rst_l(rst_l),
		.clk(busclk),
		.clken(bus_ifu_bus_clk_en),
		.rawclk(clk),
		.din(ifu_axi_rid[pt[826-:8] - 1:0]),
		.dout(ifu_bus_rid_ff[pt[826-:8] - 1:0])
	);
	rvdffe #(.WIDTH(64)) bus_data_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(clk),
		.din(ifu_axi_rdata[63:0]),
		.dout(ifu_bus_rdata_ff[63:0]),
		.en(ifu_bus_clk_en & ifu_axi_rvalid)
	);
	assign ifu_bus_cmd_ready = ifu_axi_arready;
	assign ifu_bus_rsp_valid = ifu_axi_rvalid;
	assign ifu_bus_rsp_ready = ifu_axi_rready;
	assign ifu_bus_rsp_tag[pt[826-:8] - 1:0] = ifu_axi_rid[pt[826-:8] - 1:0];
	assign ifu_bus_rsp_rdata[63:0] = ifu_axi_rdata[63:0];
	assign ifu_bus_rsp_opc[1:0] = {ifu_axi_rresp[1:0]};
	assign ifu_bus_rvalid = ifu_bus_rsp_valid & bus_ifu_bus_clk_en;
	assign ifu_bus_arready = ifu_bus_arready_unq & bus_ifu_bus_clk_en;
	assign ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff;
	assign ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff;
	assign bus_cmd_sent = ((ifu_bus_arvalid & ifu_bus_arready) & miss_pending) & ~dec_tlu_force_halt;
	assign bus_inc_data_beat_cnt = (bus_ifu_wr_en_ff & ~bus_last_data_beat) & ~dec_tlu_force_halt;
	assign bus_reset_data_beat_cnt = (ic_act_miss_f | (bus_ifu_wr_en_ff & bus_last_data_beat)) | dec_tlu_force_halt;
	assign bus_hold_data_beat_cnt = ~bus_inc_data_beat_cnt & ~bus_reset_data_beat_cnt;
	function automatic signed [pt[1174-:8] - 1:0] sv2v_cast_4BA5C_signed;
		input reg signed [pt[1174-:8] - 1:0] inp;
		sv2v_cast_4BA5C_signed = inp;
	endfunction
	assign bus_new_data_beat_count[pt[1174-:8] - 1:0] = (({pt[1174-:8] {bus_reset_data_beat_cnt}} & sv2v_cast_4BA5C_signed(0)) | ({pt[1174-:8] {bus_inc_data_beat_cnt}} & (bus_data_beat_count[pt[1174-:8] - 1:0] + {{pt[1174-:8] - 1 {1'b0}}, 1'b1}))) | ({pt[1174-:8] {bus_hold_data_beat_cnt}} & bus_data_beat_count[pt[1174-:8] - 1:0]);
	assign last_data_recieved_in = ((bus_ifu_wr_en_ff & bus_last_data_beat) & ~scnd_miss_req) | (last_data_recieved_ff & ~ic_act_miss_f);
	assign bus_new_rd_addr_count[pt[1174-:8] - 1:0] = (~miss_pending ? imb_ff[pt[1182-:8]:3] : (scnd_miss_req_q ? imb_scnd_ff[pt[1182-:8]:3] : (bus_cmd_sent ? bus_rd_addr_count[pt[1174-:8] - 1:0] + 3'b001 : bus_rd_addr_count[pt[1174-:8] - 1:0])));
	rvdff_fpga #(.WIDTH(pt[1174-:8])) bus_rd_addr_ff(
		.rst_l(rst_l),
		.clk(busclk_reset),
		.clken((bus_ifu_bus_clk_en | ic_act_miss_f) | dec_tlu_force_halt),
		.rawclk(clk),
		.din({bus_new_rd_addr_count[pt[1174-:8] - 1:0]}),
		.dout({bus_rd_addr_count[pt[1174-:8] - 1:0]})
	);
	assign bus_inc_cmd_beat_cnt = ((ifu_bus_cmd_valid & ifu_bus_cmd_ready) & miss_pending) & ~dec_tlu_force_halt;
	assign bus_reset_cmd_beat_cnt_0 = (ic_act_miss_f & ~uncacheable_miss_in) | dec_tlu_force_halt;
	assign bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in;
	assign bus_hold_cmd_beat_cnt = ~bus_inc_cmd_beat_cnt & ~((ic_act_miss_f | scnd_miss_req) | dec_tlu_force_halt);
	assign bus_cmd_beat_en = (bus_inc_cmd_beat_cnt | ic_act_miss_f) | dec_tlu_force_halt;
	function automatic [pt[1174-:8] - 1:0] sv2v_cast_4BA5C;
		input reg [pt[1174-:8] - 1:0] inp;
		sv2v_cast_4BA5C = inp;
	endfunction
	assign bus_new_cmd_beat_count[pt[1174-:8] - 1:0] = ((({pt[1174-:8] {bus_reset_cmd_beat_cnt_0}} & sv2v_cast_4BA5C_signed(0)) | ({pt[1174-:8] {bus_reset_cmd_beat_cnt_secondlast}} & sv2v_cast_4BA5C(pt[1048-:8]))) | ({pt[1174-:8] {bus_inc_cmd_beat_cnt}} & (bus_cmd_beat_count[pt[1174-:8] - 1:0] + {{pt[1174-:8] - 1 {1'b0}}, 1'b1}))) | ({pt[1174-:8] {bus_hold_cmd_beat_cnt}} & bus_cmd_beat_count[pt[1174-:8] - 1:0]);
	rvclkhdr bus_clk_reset(
		.en((bus_ifu_bus_clk_en | ic_act_miss_f) | dec_tlu_force_halt),
		.l1clk(busclk_reset),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvdffs_fpga #(.WIDTH(pt[1174-:8])) bus_cmd_beat_ff(
		.rst_l(rst_l),
		.clk(busclk_reset),
		.clken((bus_ifu_bus_clk_en | ic_act_miss_f) | dec_tlu_force_halt),
		.rawclk(clk),
		.en(bus_cmd_beat_en),
		.din({bus_new_cmd_beat_count[pt[1174-:8] - 1:0]}),
		.dout({bus_cmd_beat_count[pt[1174-:8] - 1:0]})
	);
	assign bus_last_data_beat = (uncacheable_miss_ff ? bus_data_beat_count[pt[1174-:8] - 1:0] == {{pt[1174-:8] - 1 {1'b0}}, 1'b1} : &bus_data_beat_count[pt[1174-:8] - 1:0]);
	assign bus_ifu_wr_en = ifu_bus_rvalid & miss_pending;
	assign bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending;
	assign bus_ifu_wr_en_ff_q = (((ifu_bus_rvalid_ff & miss_pending) & ~uncacheable_miss_ff) & ~(|ifu_bus_rresp_ff[1:0])) & write_ic_16_bytes;
	assign bus_ifu_wr_en_ff_wo_err = (ifu_bus_rvalid_ff & miss_pending) & ~uncacheable_miss_ff;
	rvdffie #(.WIDTH(10)) misc_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({ic_act_miss_f, ifu_wr_cumulative_err, exu_flush_final, ic_crit_wd_rdy_new_in, bus_ifu_bus_clk_en, scnd_miss_req_in, bus_cmd_req_in, last_data_recieved_in, ifc_dma_access_ok_d, dma_iccm_req}),
		.dout({ic_act_miss_f_delayed, ifu_wr_data_comb_err_ff, flush_final_f, ic_crit_wd_rdy_new_ff, bus_ifu_bus_clk_en_ff, scnd_miss_req_q, bus_cmd_req_hold, last_data_recieved_ff, ifc_dma_access_ok_prev, dma_iccm_req_f})
	);
	rvdffie #(
		.WIDTH(pt[1174-:8] + 5),
		.OVERRIDE(1)
	) misc1_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({reset_ic_in, sel_mb_addr, bus_new_data_beat_count[pt[1174-:8] - 1:0], ifc_region_acc_fault_memory_bf, ic_debug_rd_en, ic_debug_rd_en_ff}),
		.dout({reset_ic_ff, sel_mb_addr_ff, bus_data_beat_count[pt[1174-:8] - 1:0], ifc_region_acc_fault_memory_f, ic_debug_rd_en_ff, ifu_ic_debug_rd_data_valid})
	);
	assign reset_tag_valid_for_miss = (ic_act_miss_f_delayed & (miss_state == CRIT_BYP_OK)) & ~uncacheable_miss_ff;
	assign bus_ifu_wr_data_error = (|ifu_bus_rsp_opc[1:0] & ifu_bus_rvalid) & miss_pending;
	assign bus_ifu_wr_data_error_ff = (|ifu_bus_rresp_ff[1:0] & ifu_bus_rvalid_ff) & miss_pending;
	assign ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff;
	assign last_beat = bus_last_data_beat & bus_ifu_wr_en_ff;
	assign reset_beat_cnt = bus_reset_data_beat_cnt;
	assign ifc_dma_access_ok_d = (ifc_dma_access_ok & ~iccm_correct_ecc) & ~iccm_dma_sb_error;
	assign ifc_dma_access_q_ok = (((ifc_dma_access_ok & ~iccm_correct_ecc) & ifc_dma_access_ok_prev) & (perr_state == ERR_IDLE)) & ~iccm_dma_sb_error;
	assign iccm_ready = ifc_dma_access_q_ok;
	wire [1:0] iccm_ecc_word_enable;
	generate
		if (pt[927-:5] == 1) begin : iccm_enabled
			wire [3:2] dma_mem_addr_ff;
			wire iccm_dma_rden;
			wire iccm_dma_ecc_error_in;
			wire [13:0] dma_mem_ecc;
			wire [63:0] iccm_dma_rdata_in;
			wire [31:0] iccm_dma_rdata_1_muxed;
			wire [63:0] iccm_corrected_data;
			wire [13:0] iccm_corrected_ecc;
			wire [1:0] iccm_double_ecc_error;
			wire [pt[936-:9] - 1:2] iccm_rw_addr_f;
			wire [31:0] iccm_corrected_data_f_mux;
			wire [6:0] iccm_corrected_ecc_f_mux;
			wire iccm_dma_rvalid_in;
			wire [77:0] iccm_rdmux_data;
			wire iccm_rd_ecc_single_err_hold_in;
			wire [2:0] dma_mem_tag_ff;
			assign iccm_wren = ((ifc_dma_access_q_ok & dma_iccm_req) & dma_mem_write) | iccm_correct_ecc;
			assign iccm_rden = ((ifc_dma_access_q_ok & dma_iccm_req) & ~dma_mem_write) | (ifc_iccm_access_bf & ifc_fetch_req_bf);
			assign iccm_dma_rden = (ifc_dma_access_q_ok & dma_iccm_req) & ~dma_mem_write;
			assign iccm_wr_size[2:0] = {3 {dma_iccm_req}} & dma_mem_sz[2:0];
			rvecc_encode iccm_ecc_encode0(
				.din(dma_mem_wdata[31:0]),
				.ecc_out(dma_mem_ecc[6:0])
			);
			rvecc_encode iccm_ecc_encode1(
				.din(dma_mem_wdata[63:32]),
				.ecc_out(dma_mem_ecc[13:7])
			);
			assign iccm_wr_data[77:0] = (iccm_correct_ecc & ~(ifc_dma_access_q_ok & dma_iccm_req) ? {iccm_ecc_corr_data_ff[38:0], iccm_ecc_corr_data_ff[38:0]} : {dma_mem_ecc[13:7], dma_mem_wdata[63:32], dma_mem_ecc[6:0], dma_mem_wdata[31:0]});
			assign iccm_dma_rdata_1_muxed[31:0] = (dma_mem_addr_ff[2] ? iccm_corrected_data[31-:32] : iccm_corrected_data[63-:32]);
			assign iccm_dma_rdata_in[63:0] = (iccm_dma_ecc_error_in ? {2 {dma_mem_addr[31:0]}} : {iccm_dma_rdata_1_muxed[31:0], iccm_corrected_data[0+:32]});
			assign iccm_dma_ecc_error_in = |iccm_double_ecc_error[1:0];
			rvdffe #(.WIDTH(64)) dma_data_ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(clk),
				.en(iccm_dma_rvalid_in),
				.din(iccm_dma_rdata_in[63:0]),
				.dout(iccm_dma_rdata[63:0])
			);
			rvdffie #(.WIDTH(11)) dma_misc_bits(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(free_l2clk),
				.din({dma_mem_tag[2:0], dma_mem_tag_ff[2:0], dma_mem_addr[3:2], iccm_dma_rden, iccm_dma_rvalid_in, iccm_dma_ecc_error_in}),
				.dout({dma_mem_tag_ff[2:0], iccm_dma_rtag[2:0], dma_mem_addr_ff[3:2], iccm_dma_rvalid_in, iccm_dma_rvalid, iccm_dma_ecc_error})
			);
			assign iccm_rw_addr[pt[936-:9] - 1:1] = ((ifc_dma_access_q_ok & dma_iccm_req) & ~iccm_correct_ecc ? dma_mem_addr[pt[936-:9] - 1:1] : (~(ifc_dma_access_q_ok & dma_iccm_req) & iccm_correct_ecc ? {iccm_ecc_corr_index_ff[pt[936-:9] - 1:2], 1'b0} : ifc_fetch_addr_bf[pt[936-:9] - 1:1]));
			wire [3:0] ic_fetch_val_int_f;
			wire [3:0] ic_fetch_val_shift_right;
			assign ic_fetch_val_int_f[3:0] = {2'b00, ic_fetch_val_f[1:0]};
			assign ic_fetch_val_shift_right[3:0] = {ic_fetch_val_int_f << ifu_fetch_addr_int_f[1]};
			assign iccm_rdmux_data[77:0] = iccm_rd_data_ecc[77:0];
			for (i = 0; i < 2; i = i + 1) begin : ICCM_ECC_CHECK
				assign iccm_ecc_word_enable[i] = (((|ic_fetch_val_shift_right[(2 * i) + 1:2 * i] & ~exu_flush_final) & sel_iccm_data) | iccm_dma_rvalid_in) & ~dec_tlu_core_ecc_disable;
				rvecc_decode ecc_decode(
					.en(iccm_ecc_word_enable[i]),
					.sed_ded(1'b0),
					.din(iccm_rdmux_data[(39 * i) + 31:39 * i]),
					.ecc_in(iccm_rdmux_data[(39 * i) + 38:(39 * i) + 32]),
					.dout(iccm_corrected_data[(i * 32) + 31-:32]),
					.ecc_out(iccm_corrected_ecc[(i * 7) + 6-:7]),
					.single_ecc_error(iccm_single_ecc_error[i]),
					.double_ecc_error(iccm_double_ecc_error[i])
				);
			end
			assign iccm_rd_ecc_single_err = (|iccm_single_ecc_error[1:0] & ifc_iccm_access_f) & ifc_fetch_req_f;
			assign iccm_rd_ecc_double_err[1:0] = (~ifu_fetch_addr_int_f[1] ? {iccm_double_ecc_error[0], iccm_double_ecc_error[0]} & {2 {ifc_iccm_access_f}} : {iccm_double_ecc_error[1], iccm_double_ecc_error[0]} & {2 {ifc_iccm_access_f}});
			assign iccm_corrected_data_f_mux[31:0] = (iccm_single_ecc_error[0] ? iccm_corrected_data[0+:32] : iccm_corrected_data[32+:32]);
			assign iccm_corrected_ecc_f_mux[6:0] = (iccm_single_ecc_error[0] ? iccm_corrected_ecc[0+:7] : iccm_corrected_ecc[7+:7]);
			assign iccm_ecc_write_status = ((iccm_rd_ecc_single_err & ~iccm_rd_ecc_single_err_ff) & ~exu_flush_final) | iccm_dma_sb_error;
			assign iccm_rd_ecc_single_err_hold_in = (iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff) & ~exu_flush_final;
			assign iccm_error_start = iccm_rd_ecc_single_err;
			assign iccm_ecc_corr_index_in[pt[936-:9] - 1:2] = (iccm_single_ecc_error[0] ? iccm_rw_addr_f[pt[936-:9] - 1:2] : iccm_rw_addr_f[pt[936-:9] - 1:2] + 1'b1);
			rvdffie #(.WIDTH(pt[936-:9] - 1)) iccm_index_f(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(free_l2clk),
				.din({iccm_rw_addr[pt[936-:9] - 1:2], iccm_rd_ecc_single_err_hold_in}),
				.dout({iccm_rw_addr_f[pt[936-:9] - 1:2], iccm_rd_ecc_single_err_ff})
			);
			rvdffe #(.WIDTH(pt[936-:9] + 37)) ecc_dat0_ff(
				.clk(clk),
				.din({iccm_corrected_ecc_f_mux[6:0], iccm_corrected_data_f_mux[31:0], iccm_ecc_corr_index_in[pt[936-:9] - 1:2]}),
				.dout({iccm_ecc_corr_data_ff[38:0], iccm_ecc_corr_index_ff[pt[936-:9] - 1:2]}),
				.en(iccm_ecc_write_status),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
		end
		else begin : iccm_disabled
			assign iccm_dma_rvalid = 1'b0;
			assign iccm_dma_ecc_error = 1'b0;
			assign iccm_dma_rdata[63:0] = {64 {1'sb0}};
			assign iccm_single_ecc_error = {2 {1'sb0}};
			assign iccm_dma_rtag = {3 {1'sb0}};
			assign iccm_rd_ecc_single_err = 1'b0;
			assign iccm_rd_ecc_double_err = {2 {1'sb0}};
			assign iccm_rd_ecc_single_err_ff = 1'b0;
			assign iccm_error_start = 1'b0;
			assign iccm_ecc_corr_index_ff[pt[936-:9] - 1:2] = {((pt[936-:9] - 1) >= 2 ? pt[936-:9] - 2 : 4 - pt[936-:9]) {1'sb0}};
			assign iccm_ecc_corr_data_ff[38:0] = {39 {1'sb0}};
			assign iccm_ecc_write_status = 1'b0;
		end
	endgenerate
	assign ic_rd_en = (((ifc_fetch_req_bf & ~ifc_fetch_uncacheable_bf) & ~ifc_iccm_access_bf) & ~(((((((miss_state == STREAM) & ~miss_state_en) | ((miss_state == CRIT_BYP_OK) & ~miss_state_en)) | ((miss_state == STALL_SCND_MISS) & ~miss_state_en)) | ((miss_state == MISS_WAIT) & ~miss_state_en)) | ((miss_state == CRIT_WRD_RDY) & ~miss_state_en)) | (((miss_state == CRIT_BYP_OK) & miss_state_en) & (miss_nxtstate == MISS_WAIT)))) | (((ifc_fetch_req_bf & exu_flush_final) & ~ifc_fetch_uncacheable_bf) & ~ifc_iccm_access_bf);
	wire ic_real_rd_wp_unused;
	assign ic_real_rd_wp_unused = ((((((ifc_fetch_req_bf & ~ifc_iccm_access_bf) & ~ifc_region_acc_fault_final_bf) & ~dec_tlu_fence_i_wb) & ~stream_miss_f) & ~ic_act_miss_f) & ~(((((((((miss_state == STREAM) & ~miss_state_en) | (((miss_state == CRIT_BYP_OK) & ~miss_state_en) & ~(miss_nxtstate == MISS_WAIT))) | (((miss_state == CRIT_BYP_OK) & miss_state_en) & (miss_nxtstate == MISS_WAIT))) | ((miss_state == MISS_WAIT) & ~miss_state_en)) | ((miss_state == STALL_SCND_MISS) & ~miss_state_en)) | ((miss_state == CRIT_WRD_RDY) & ~miss_state_en)) | ((miss_nxtstate == STREAM) & miss_state_en)) | ((miss_state == SCND_MISS) & ~miss_state_en))) | (((((ifc_fetch_req_bf & ~ifc_iccm_access_bf) & ~ifc_region_acc_fault_final_bf) & ~dec_tlu_fence_i_wb) & ~stream_miss_f) & exu_flush_final);
	assign ic_wr_en[pt[1060-:7] - 1:0] = bus_ic_wr_en[pt[1060-:7] - 1:0] & {pt[1060-:7] {write_ic_16_bytes}};
	assign ic_write_stall = write_ic_16_bytes & ~(((miss_state == CRIT_BYP_OK) | ((miss_state == STREAM) & ~((exu_flush_final | ifu_bp_hit_taken_q_f) | stream_eol_f))) & ~((bus_ifu_wr_en_ff & last_beat) & ~uncacheable_miss_ff));
	reg [pt[1060-:7] - 1:0] ic_tag_valid_unq;
	generate
		if (pt[1120-:5] == 1) begin : icache_enabled
			assign ic_valid = (~ifu_wr_cumulative_err_data & ~(reset_ic_in | reset_ic_ff)) & ~reset_tag_valid_for_miss;
			assign ifu_status_wr_addr_w_debug[pt[1104-:9]:pt[998-:7]] = ((ic_debug_rd_en | ic_debug_wr_en) & ic_debug_tag_array ? ic_debug_addr[pt[1104-:9]:pt[998-:7]] : ifu_status_wr_addr[pt[1104-:9]:pt[998-:7]]);
			assign way_status_wr_en_w_debug = way_status_wr_en | (ic_debug_wr_en & ic_debug_tag_array);
			assign way_status_new_w_debug[pt[1027-:7] - 1:0] = (ic_debug_wr_en & ic_debug_tag_array ? (pt[1027-:7] == 1 ? ic_debug_wr_data[4] : ic_debug_wr_data[6:4]) : way_status_new[pt[1027-:7] - 1:0]);
			rvdffie #(
				.WIDTH(((pt[991-:9] - pt[998-:7]) + 1) + pt[1027-:7]),
				.OVERRIDE(1)
			) status_misc_ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(free_l2clk),
				.din({ifu_status_wr_addr_w_debug[pt[1104-:9]:pt[998-:7]], way_status_wr_en_w_debug, way_status_new_w_debug[pt[1027-:7] - 1:0]}),
				.dout({ifu_status_wr_addr_ff[pt[1104-:9]:pt[998-:7]], way_status_wr_en_ff, way_status_new_ff[pt[1027-:7] - 1:0]})
			);
			wire [(pt[1015-:17] / 8) - 1:0] way_status_clken;
			wire [(pt[1015-:17] / 8) - 1:0] way_status_clk;
			for (i = 0; i < (pt[1015-:17] / 8); i = i + 1) begin : CLK_GRP_WAY_STATUS
				assign way_status_clken[i] = ifu_status_wr_addr_ff[pt[1104-:9]:pt[998-:7] + 3] == i;
				rvclkhdr way_status_cgc(
					.en(way_status_clken[i]),
					.l1clk(way_status_clk[i]),
					.clk(clk),
					.scan_mode(scan_mode)
				);
				genvar j;
				for (j = 0; j < 8; j = j + 1) begin : WAY_STATUS
					rvdffs_fpga #(.WIDTH(pt[1027-:7])) ic_way_status(
						.rst_l(rst_l),
						.clk(way_status_clk[i]),
						.clken(way_status_clken[i]),
						.rawclk(clk),
						.en((ifu_status_wr_addr_ff[pt[998-:7] + 2:pt[998-:7]] == j) & way_status_wr_en_ff),
						.din(way_status_new_ff[pt[1027-:7] - 1:0]),
						.dout(way_status_out[((8 * i) + j) * pt[1027-:7]+:pt[1027-:7]])
					);
				end
			end
			function automatic signed [(pt[991-:9] - pt[998-:7]) - 1:0] sv2v_cast_46E4F_signed;
				input reg signed [(pt[991-:9] - pt[998-:7]) - 1:0] inp;
				sv2v_cast_46E4F_signed = inp;
			endfunction
			always @(*) begin : way_status_out_mux
				way_status[pt[1027-:7] - 1:0] = {pt[1027-:7] {1'sb0}};
				begin : sv2v_autoblock_47
					reg signed [31:0] j;
					for (j = 0; j < pt[1015-:17]; j = j + 1)
						begin : status_mux_loop
							if (ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7]] == sv2v_cast_46E4F_signed(j)) begin : mux_out
								way_status[pt[1027-:7] - 1:0] = way_status_out[j * pt[1027-:7]+:pt[1027-:7]];
							end
						end
				end
			end
			assign ifu_ic_rw_int_addr_w_debug[pt[1104-:9]:pt[998-:7]] = ((ic_debug_rd_en | ic_debug_wr_en) & ic_debug_tag_array ? ic_debug_addr[pt[1104-:9]:pt[998-:7]] : ifu_ic_rw_int_addr[pt[1104-:9]:pt[998-:7]]);
			assign ifu_tag_wren_w_debug[pt[1060-:7] - 1:0] = ifu_tag_wren[pt[1060-:7] - 1:0] | ic_debug_tag_wr_en[pt[1060-:7] - 1:0];
			assign ic_valid_w_debug = (ic_debug_wr_en & ic_debug_tag_array ? ic_debug_wr_data[0] : ic_valid);
			rvdffie #(.WIDTH(((pt[991-:9] - pt[998-:7]) + pt[1060-:7]) + 1)) tag_addr_ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.clk(free_l2clk),
				.din({ifu_ic_rw_int_addr_w_debug[pt[1104-:9]:pt[998-:7]], ifu_tag_wren_w_debug[pt[1060-:7] - 1:0], ic_valid_w_debug}),
				.dout({ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7]], ifu_tag_wren_ff[pt[1060-:7] - 1:0], ic_valid_ff})
			);
			wire [(pt[1060-:7] * pt[1015-:17]) - 1:0] ic_tag_valid_out;
			wire [((pt[1015-:17] / 32) * pt[1060-:7]) - 1:0] tag_valid_clken;
			wire [((pt[1015-:17] / 32) * pt[1060-:7]) - 1:0] tag_valid_clk;
			for (i = 0; i < (pt[1015-:17] / 32); i = i + 1) begin : CLK_GRP_TAG_VALID
				genvar j;
				for (j = 0; j < pt[1060-:7]; j = j + 1) begin : way_clken
					if (pt[1015-:17] == 32) begin
						assign tag_valid_clken[(i * pt[1060-:7]) + j] = (ifu_tag_wren_ff[j] | perr_err_inv_way[j]) | reset_all_tags;
					end
					else assign tag_valid_clken[(i * pt[1060-:7]) + j] = (((ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7] + 5] == i) & ifu_tag_wren_ff[j]) | ((perr_ic_index_ff[pt[1104-:9]:pt[998-:7] + 5] == i) & perr_err_inv_way[j])) | reset_all_tags;
					rvclkhdr way_status_cgc(
						.en(tag_valid_clken[(i * pt[1060-:7]) + j]),
						.l1clk(tag_valid_clk[(i * pt[1060-:7]) + j]),
						.clk(clk),
						.scan_mode(scan_mode)
					);
					genvar k;
					for (k = 0; k < 32; k = k + 1) begin : TAG_VALID
						rvdffs_fpga #(.WIDTH(1)) ic_way_tagvalid_dup(
							.rst_l(rst_l),
							.clk(tag_valid_clk[(i * pt[1060-:7]) + j]),
							.clken(tag_valid_clken[(i * pt[1060-:7]) + j]),
							.rawclk(clk),
							.en((((ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7]] == (k + (32 * i))) & ifu_tag_wren_ff[j]) | ((perr_ic_index_ff[pt[1104-:9]:pt[998-:7]] == (k + (32 * i))) & perr_err_inv_way[j])) | reset_all_tags),
							.din((ic_valid_ff & ~reset_all_tags) & ~perr_sel_invalidate),
							.dout(ic_tag_valid_out[(j * pt[1015-:17]) + ((32 * i) + k)])
						);
					end
				end
			end
			always @(*) begin : tag_valid_out_mux
				ic_tag_valid_unq[pt[1060-:7] - 1:0] = {pt[1060-:7] {1'sb0}};
				begin : sv2v_autoblock_48
					reg signed [31:0] j;
					for (j = 0; j < pt[1015-:17]; j = j + 1)
						begin : tag_valid_loop
							if (ifu_ic_rw_int_addr_ff[pt[1104-:9]:pt[998-:7]] == sv2v_cast_46E4F_signed(j)) begin : valid_out
								begin : sv2v_autoblock_49
									reg signed [31:0] k;
									for (k = 0; k < pt[1060-:7]; k = k + 1)
										ic_tag_valid_unq[k] = ic_tag_valid_unq[k] | ic_tag_valid_out[(k * pt[1015-:17]) + j];
								end
							end
						end
				end
			end
			if (pt[1060-:7] == 4) begin : four_way_plru
				assign replace_way_mb_any[3] = ((way_status_mb_ff[2] & way_status_mb_ff[0]) & &tagv_mb_ff[3:0]) | (((~tagv_mb_ff[3] & tagv_mb_ff[2]) & tagv_mb_ff[1]) & tagv_mb_ff[0]);
				assign replace_way_mb_any[2] = ((~way_status_mb_ff[2] & way_status_mb_ff[0]) & &tagv_mb_ff[3:0]) | ((~tagv_mb_ff[2] & tagv_mb_ff[1]) & tagv_mb_ff[0]);
				assign replace_way_mb_any[1] = ((way_status_mb_ff[1] & ~way_status_mb_ff[0]) & &tagv_mb_ff[3:0]) | (~tagv_mb_ff[1] & tagv_mb_ff[0]);
				assign replace_way_mb_any[0] = ((~way_status_mb_ff[1] & ~way_status_mb_ff[0]) & &tagv_mb_ff[3:0]) | ~tagv_mb_ff[0];
				assign way_status_hit_new[pt[1027-:7] - 1:0] = ((({3 {~exu_flush_final & ic_rd_hit[0]}} & {way_status[2], 1'b1, 1'b1}) | ({3 {~exu_flush_final & ic_rd_hit[1]}} & {way_status[2], 1'b0, 1'b1})) | ({3 {~exu_flush_final & ic_rd_hit[2]}} & {1'b1, way_status[1], 1'b0})) | ({3 {~exu_flush_final & ic_rd_hit[3]}} & {1'b0, way_status[1], 1'b0});
				assign way_status_rep_new[pt[1027-:7] - 1:0] = ((({3 {replace_way_mb_any[0]}} & {way_status_mb_ff[2], 1'b1, 1'b1}) | ({3 {replace_way_mb_any[1]}} & {way_status_mb_ff[2], 1'b0, 1'b1})) | ({3 {replace_way_mb_any[2]}} & {1'b1, way_status_mb_ff[1], 1'b0})) | ({3 {replace_way_mb_any[3]}} & {1'b0, way_status_mb_ff[1], 1'b0});
			end
			else begin : two_ways_plru
				assign replace_way_mb_any[0] = ((~way_status_mb_ff & tagv_mb_ff[0]) & tagv_mb_ff[1]) | ~tagv_mb_ff[0];
				assign replace_way_mb_any[1] = ((way_status_mb_ff & tagv_mb_ff[0]) & tagv_mb_ff[1]) | (~tagv_mb_ff[1] & tagv_mb_ff[0]);
				assign way_status_hit_new[pt[1027-:7] - 1:0] = ic_rd_hit[0];
				assign way_status_rep_new[pt[1027-:7] - 1:0] = replace_way_mb_any[0];
			end
			assign way_status_new[pt[1027-:7] - 1:0] = (bus_ifu_wr_en_ff_q & last_beat ? way_status_rep_new[pt[1027-:7] - 1:0] : way_status_hit_new[pt[1027-:7] - 1:0]);
			assign way_status_wr_en = (bus_ifu_wr_en_ff_q & last_beat) | ic_act_hit_f;
			for (i = 0; i < pt[1060-:7]; i = i + 1) begin : bus_wren_loop
				assign bus_wren[i] = (bus_ifu_wr_en_ff_q & replace_way_mb_any[i]) & miss_pending;
				assign bus_wren_last[i] = ((bus_ifu_wr_en_ff_wo_err & replace_way_mb_any[i]) & miss_pending) & bus_last_data_beat;
				assign ifu_tag_wren[i] = bus_wren_last[i] | wren_reset_miss[i];
				assign wren_reset_miss[i] = replace_way_mb_any[i] & reset_tag_valid_for_miss;
			end
			assign bus_ic_wr_en[pt[1060-:7] - 1:0] = bus_wren[pt[1060-:7] - 1:0];
		end
		else begin : icache_disabled
			wire [pt[1060-:7]:1] sv2v_tmp_602A9;
			assign sv2v_tmp_602A9 = {pt[1060-:7] {1'sb0}};
			always @(*) ic_tag_valid_unq[pt[1060-:7] - 1:0] = sv2v_tmp_602A9;
			wire [pt[1027-:7]:1] sv2v_tmp_89B17;
			assign sv2v_tmp_89B17 = {pt[1027-:7] {1'sb0}};
			always @(*) way_status[pt[1027-:7] - 1:0] = sv2v_tmp_89B17;
			assign replace_way_mb_any[pt[1060-:7] - 1:0] = {pt[1060-:7] {1'sb0}};
			assign way_status_hit_new[pt[1027-:7] - 1:0] = {pt[1027-:7] {1'sb0}};
			assign way_status_rep_new[pt[1027-:7] - 1:0] = {pt[1027-:7] {1'sb0}};
			assign way_status_new[pt[1027-:7] - 1:0] = {pt[1027-:7] {1'sb0}};
			assign way_status_wr_en = 1'b0;
			assign bus_wren[pt[1060-:7] - 1:0] = {pt[1060-:7] {1'sb0}};
		end
	endgenerate
	assign ic_tag_valid[pt[1060-:7] - 1:0] = ic_tag_valid_unq[pt[1060-:7] - 1:0] & {pt[1060-:7] {~fetch_uncacheable_ff & ifc_fetch_req_f_raw}};
	assign ic_debug_tag_val_rd_out = |((ic_tag_valid_unq[pt[1060-:7] - 1:0] & ic_debug_way_ff[pt[1060-:7] - 1:0]) & {pt[1060-:7] {ic_debug_rd_en_ff}});
	assign ifu_pmu_ic_miss_in = ic_act_miss_f;
	assign ifu_pmu_ic_hit_in = ic_act_hit_f;
	assign ifu_pmu_bus_error_in = |ifc_bus_acc_fault_f;
	assign ifu_pmu_bus_trxn_in = bus_cmd_sent;
	assign ifu_pmu_bus_busy_in = (ifu_bus_arvalid_ff & ~ifu_bus_arready_ff) & miss_pending;
	rvdffie #(.WIDTH(9)) ifu_pmu_sigs_ff(
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.clk(free_l2clk),
		.din({ifc_fetch_uncacheable_bf, ifc_fetch_req_qual_bf, dma_sb_err_state, dec_tlu_fence_i_wb, ifu_pmu_ic_miss_in, ifu_pmu_ic_hit_in, ifu_pmu_bus_error_in, ifu_pmu_bus_busy_in, ifu_pmu_bus_trxn_in}),
		.dout({fetch_uncacheable_ff, ifc_fetch_req_f_raw, dma_sb_err_state_ff, reset_all_tags, ifu_pmu_ic_miss, ifu_pmu_ic_hit, ifu_pmu_bus_error, ifu_pmu_bus_busy, ifu_pmu_bus_trxn})
	);
	assign ic_debug_addr[pt[1104-:9]:3] = dec_tlu_ic_diag_pkt[pt[1104-:9] - 1:2];
	assign ic_debug_way_enc[1:0] = dec_tlu_ic_diag_pkt[17:16];
	assign ic_debug_tag_array = dec_tlu_ic_diag_pkt[18];
	assign ic_debug_rd_en = dec_tlu_ic_diag_pkt[1];
	assign ic_debug_wr_en = dec_tlu_ic_diag_pkt[0];
	assign ic_debug_way[pt[1060-:7] - 1:0] = {ic_debug_way_enc[1:0] == 2'b11, ic_debug_way_enc[1:0] == 2'b10, ic_debug_way_enc[1:0] == 2'b01, ic_debug_way_enc[1:0] == 2'b00};
	assign ic_debug_tag_wr_en[pt[1060-:7] - 1:0] = {pt[1060-:7] {ic_debug_wr_en & ic_debug_tag_array}} & ic_debug_way[pt[1060-:7] - 1:0];
	assign ic_debug_ict_array_sel_in = ic_debug_rd_en & ic_debug_tag_array;
	rvdff_fpga #(.WIDTH(1 + pt[1060-:7])) ifu_debug_sel_ff(
		.rst_l(rst_l),
		.clk(debug_c1_clk),
		.clken(debug_c1_clken),
		.rawclk(clk),
		.din({ic_debug_ict_array_sel_in, ic_debug_way[pt[1060-:7] - 1:0]}),
		.dout({ic_debug_ict_array_sel_ff, ic_debug_way_ff[pt[1060-:7] - 1:0]})
	);
	assign debug_data_clken = ic_debug_rd_en_ff;
	assign ifc_region_acc_okay = (((((((~(|{pt[530-:5], pt[525-:5], pt[520-:5], pt[515-:5], pt[510-:5], pt[505-:5], pt[500-:5], pt[495-:5]}) | (pt[530-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[490-:36]) == (pt[818-:36] | pt[490-:36])))) | (pt[525-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[454-:36]) == (pt[782-:36] | pt[454-:36])))) | (pt[520-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[418-:36]) == (pt[746-:36] | pt[418-:36])))) | (pt[515-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[382-:36]) == (pt[710-:36] | pt[382-:36])))) | (pt[510-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[346-:36]) == (pt[674-:36] | pt[346-:36])))) | (pt[505-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[310-:36]) == (pt[638-:36] | pt[310-:36])))) | (pt[500-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[274-:36]) == (pt[602-:36] | pt[274-:36])))) | (pt[495-:5] & (({ifc_fetch_addr_bf[31:1], 1'b0} | pt[238-:36]) == (pt[566-:36] | pt[238-:36])));
	assign ifc_region_acc_fault_memory_bf = (~ifc_iccm_access_bf & ~ifc_region_acc_okay) & ifc_fetch_req_bf;
	assign ifc_region_acc_fault_final_bf = ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
endmodule
module eb1_lsu (
	clk_override,
	dec_tlu_flush_lower_r,
	dec_tlu_i0_kill_writeb_r,
	dec_tlu_force_halt,
	dec_tlu_external_ldfwd_disable,
	dec_tlu_wb_coalescing_disable,
	dec_tlu_sideeffect_posted_disable,
	dec_tlu_core_ecc_disable,
	exu_lsu_rs1_d,
	exu_lsu_rs2_d,
	dec_lsu_offset_d,
	lsu_p,
	dec_lsu_valid_raw_d,
	dec_tlu_mrac_ff,
	lsu_result_m,
	lsu_result_corr_r,
	lsu_load_stall_any,
	lsu_store_stall_any,
	lsu_fastint_stall_any,
	lsu_idle_any,
	lsu_active,
	lsu_fir_addr,
	lsu_fir_error,
	lsu_single_ecc_error_incr,
	lsu_error_pkt_r,
	lsu_imprecise_error_load_any,
	lsu_imprecise_error_store_any,
	lsu_imprecise_error_addr_any,
	lsu_nonblock_load_valid_m,
	lsu_nonblock_load_tag_m,
	lsu_nonblock_load_inv_r,
	lsu_nonblock_load_inv_tag_r,
	lsu_nonblock_load_data_valid,
	lsu_nonblock_load_data_error,
	lsu_nonblock_load_data_tag,
	lsu_nonblock_load_data,
	lsu_pmu_load_external_m,
	lsu_pmu_store_external_m,
	lsu_pmu_misaligned_m,
	lsu_pmu_bus_trxn,
	lsu_pmu_bus_misaligned,
	lsu_pmu_bus_error,
	lsu_pmu_bus_busy,
	trigger_pkt_any,
	lsu_trigger_match_m,
	dccm_wren,
	dccm_rden,
	dccm_wr_addr_lo,
	dccm_wr_addr_hi,
	dccm_rd_addr_lo,
	dccm_rd_addr_hi,
	dccm_wr_data_lo,
	dccm_wr_data_hi,
	dccm_rd_data_lo,
	dccm_rd_data_hi,
	picm_wren,
	picm_rden,
	picm_mken,
	picm_rdaddr,
	picm_wraddr,
	picm_wr_data,
	picm_rd_data,
	lsu_axi_awvalid,
	lsu_axi_awready,
	lsu_axi_awid,
	lsu_axi_awaddr,
	lsu_axi_awregion,
	lsu_axi_awlen,
	lsu_axi_awsize,
	lsu_axi_awburst,
	lsu_axi_awlock,
	lsu_axi_awcache,
	lsu_axi_awprot,
	lsu_axi_awqos,
	lsu_axi_wvalid,
	lsu_axi_wready,
	lsu_axi_wdata,
	lsu_axi_wstrb,
	lsu_axi_wlast,
	lsu_axi_bvalid,
	lsu_axi_bready,
	lsu_axi_bresp,
	lsu_axi_bid,
	lsu_axi_arvalid,
	lsu_axi_arready,
	lsu_axi_arid,
	lsu_axi_araddr,
	lsu_axi_arregion,
	lsu_axi_arlen,
	lsu_axi_arsize,
	lsu_axi_arburst,
	lsu_axi_arlock,
	lsu_axi_arcache,
	lsu_axi_arprot,
	lsu_axi_arqos,
	lsu_axi_rvalid,
	lsu_axi_rready,
	lsu_axi_rid,
	lsu_axi_rdata,
	lsu_axi_rresp,
	lsu_axi_rlast,
	lsu_bus_clk_en,
	dma_dccm_req,
	dma_mem_tag,
	dma_mem_addr,
	dma_mem_sz,
	dma_mem_write,
	dma_mem_wdata,
	dccm_dma_rvalid,
	dccm_dma_ecc_error,
	dccm_dma_rtag,
	dccm_dma_rdata,
	dccm_ready,
	scan_mode,
	clk,
	active_clk,
	rst_l
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk_override;
	input wire dec_tlu_flush_lower_r;
	input wire dec_tlu_i0_kill_writeb_r;
	input wire dec_tlu_force_halt;
	input wire dec_tlu_external_ldfwd_disable;
	input wire dec_tlu_wb_coalescing_disable;
	input wire dec_tlu_sideeffect_posted_disable;
	input wire dec_tlu_core_ecc_disable;
	input wire [31:0] exu_lsu_rs1_d;
	input wire [31:0] exu_lsu_rs2_d;
	input wire [11:0] dec_lsu_offset_d;
	input wire [13:0] lsu_p;
	input wire dec_lsu_valid_raw_d;
	input wire [31:0] dec_tlu_mrac_ff;
	output wire [31:0] lsu_result_m;
	output wire [31:0] lsu_result_corr_r;
	output wire lsu_load_stall_any;
	output wire lsu_store_stall_any;
	output wire lsu_fastint_stall_any;
	output wire lsu_idle_any;
	output wire lsu_active;
	output wire [31:1] lsu_fir_addr;
	output wire [1:0] lsu_fir_error;
	output wire lsu_single_ecc_error_incr;
	output wire [39:0] lsu_error_pkt_r;
	output wire lsu_imprecise_error_load_any;
	output wire lsu_imprecise_error_store_any;
	output wire [31:0] lsu_imprecise_error_addr_any;
	output wire lsu_nonblock_load_valid_m;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	output wire lsu_nonblock_load_inv_r;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	output wire lsu_nonblock_load_data_valid;
	output wire lsu_nonblock_load_data_error;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	output wire [31:0] lsu_nonblock_load_data;
	output wire lsu_pmu_load_external_m;
	output wire lsu_pmu_store_external_m;
	output wire lsu_pmu_misaligned_m;
	output wire lsu_pmu_bus_trxn;
	output wire lsu_pmu_bus_misaligned;
	output wire lsu_pmu_bus_error;
	output wire lsu_pmu_bus_busy;
	input wire [151:0] trigger_pkt_any;
	output wire [3:0] lsu_trigger_match_m;
	output wire dccm_wren;
	output wire dccm_rden;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	output wire picm_wren;
	output wire picm_rden;
	output wire picm_mken;
	output wire [31:0] picm_rdaddr;
	output wire [31:0] picm_wraddr;
	output wire [31:0] picm_wr_data;
	input wire [31:0] picm_rd_data;
	output wire lsu_axi_awvalid;
	input wire lsu_axi_awready;
	output wire [pt[181-:8] - 1:0] lsu_axi_awid;
	output wire [31:0] lsu_axi_awaddr;
	output wire [3:0] lsu_axi_awregion;
	output wire [7:0] lsu_axi_awlen;
	output wire [2:0] lsu_axi_awsize;
	output wire [1:0] lsu_axi_awburst;
	output wire lsu_axi_awlock;
	output wire [3:0] lsu_axi_awcache;
	output wire [2:0] lsu_axi_awprot;
	output wire [3:0] lsu_axi_awqos;
	output wire lsu_axi_wvalid;
	input wire lsu_axi_wready;
	output wire [63:0] lsu_axi_wdata;
	output wire [7:0] lsu_axi_wstrb;
	output wire lsu_axi_wlast;
	input wire lsu_axi_bvalid;
	output wire lsu_axi_bready;
	input wire [1:0] lsu_axi_bresp;
	input wire [pt[181-:8] - 1:0] lsu_axi_bid;
	output wire lsu_axi_arvalid;
	input wire lsu_axi_arready;
	output wire [pt[181-:8] - 1:0] lsu_axi_arid;
	output wire [31:0] lsu_axi_araddr;
	output wire [3:0] lsu_axi_arregion;
	output wire [7:0] lsu_axi_arlen;
	output wire [2:0] lsu_axi_arsize;
	output wire [1:0] lsu_axi_arburst;
	output wire lsu_axi_arlock;
	output wire [3:0] lsu_axi_arcache;
	output wire [2:0] lsu_axi_arprot;
	output wire [3:0] lsu_axi_arqos;
	input wire lsu_axi_rvalid;
	output wire lsu_axi_rready;
	input wire [pt[181-:8] - 1:0] lsu_axi_rid;
	input wire [63:0] lsu_axi_rdata;
	input wire [1:0] lsu_axi_rresp;
	input wire lsu_axi_rlast;
	input wire lsu_bus_clk_en;
	input wire dma_dccm_req;
	input wire [2:0] dma_mem_tag;
	input wire [31:0] dma_mem_addr;
	input wire [2:0] dma_mem_sz;
	input wire dma_mem_write;
	input wire [63:0] dma_mem_wdata;
	output wire dccm_dma_rvalid;
	output wire dccm_dma_ecc_error;
	output wire [2:0] dccm_dma_rtag;
	output wire [63:0] dccm_dma_rdata;
	output wire dccm_ready;
	input wire scan_mode;
	input wire clk;
	input wire active_clk;
	input wire rst_l;
	wire lsu_dccm_rden_m;
	wire lsu_dccm_rden_r;
	wire [31:0] store_data_m;
	wire [31:0] store_data_r;
	wire [31:0] store_data_hi_r;
	wire [31:0] store_data_lo_r;
	wire [31:0] store_datafn_hi_r;
	wire [31:0] store_datafn_lo_r;
	wire [31:0] sec_data_lo_m;
	wire [31:0] sec_data_hi_m;
	wire [31:0] sec_data_lo_r;
	wire [31:0] sec_data_hi_r;
	wire [31:0] lsu_ld_data_m;
	wire [31:0] dccm_rdata_hi_m;
	wire [31:0] dccm_rdata_lo_m;
	wire [6:0] dccm_data_ecc_hi_m;
	wire [6:0] dccm_data_ecc_lo_m;
	wire lsu_single_ecc_error_m;
	wire lsu_double_ecc_error_m;
	wire [31:0] lsu_ld_data_r;
	wire [31:0] lsu_ld_data_corr_r;
	wire [31:0] dccm_rdata_hi_r;
	wire [31:0] dccm_rdata_lo_r;
	wire [6:0] dccm_data_ecc_hi_r;
	wire [6:0] dccm_data_ecc_lo_r;
	wire single_ecc_error_hi_r;
	wire single_ecc_error_lo_r;
	wire lsu_single_ecc_error_r;
	wire lsu_double_ecc_error_r;
	wire ld_single_ecc_error_r;
	wire ld_single_ecc_error_r_ff;
	wire [31:0] picm_mask_data_m;
	wire [31:0] lsu_addr_d;
	wire [31:0] lsu_addr_m;
	wire [31:0] lsu_addr_r;
	wire [31:0] end_addr_d;
	wire [31:0] end_addr_m;
	wire [31:0] end_addr_r;
	wire [13:0] lsu_pkt_d;
	wire [13:0] lsu_pkt_m;
	wire [13:0] lsu_pkt_r;
	wire lsu_i0_valid_d;
	wire lsu_i0_valid_m;
	wire lsu_i0_valid_r;
	wire store_stbuf_reqvld_r;
	wire ldst_stbuf_reqvld_r;
	wire lsu_commit_r;
	wire lsu_exc_m;
	wire addr_in_dccm_d;
	wire addr_in_dccm_m;
	wire addr_in_dccm_r;
	wire addr_in_pic_d;
	wire addr_in_pic_m;
	wire addr_in_pic_r;
	wire ldst_dual_d;
	wire ldst_dual_m;
	wire ldst_dual_r;
	wire addr_external_m;
	wire stbuf_reqvld_any;
	wire stbuf_reqvld_flushed_any;
	wire [pt[157-:9] - 1:0] stbuf_addr_any;
	wire [pt[1382-:10] - 1:0] stbuf_data_any;
	wire [pt[1372-:7] - 1:0] stbuf_ecc_any;
	wire [pt[1382-:10] - 1:0] sec_data_lo_r_ff;
	wire [pt[1382-:10] - 1:0] sec_data_hi_r_ff;
	wire [pt[1372-:7] - 1:0] sec_data_ecc_hi_r_ff;
	wire [pt[1372-:7] - 1:0] sec_data_ecc_lo_r_ff;
	wire lsu_cmpen_m;
	wire [pt[1382-:10] - 1:0] stbuf_fwddata_hi_m;
	wire [pt[1382-:10] - 1:0] stbuf_fwddata_lo_m;
	wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_hi_m;
	wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_lo_m;
	wire lsu_stbuf_commit_any;
	wire lsu_stbuf_empty_any;
	wire lsu_stbuf_full_any;
	wire lsu_busreq_r;
	wire lsu_bus_buffer_pend_any;
	wire lsu_bus_buffer_empty_any;
	wire lsu_bus_buffer_full_any;
	wire lsu_busreq_m;
	wire [31:0] bus_read_data_m;
	wire flush_m_up;
	wire flush_r;
	wire is_sideeffects_m;
	wire [2:0] dma_mem_tag_d;
	wire [2:0] dma_mem_tag_m;
	wire ldst_nodma_mtor;
	wire dma_dccm_wen;
	wire dma_pic_wen;
	wire [31:0] dma_dccm_wdata_lo;
	wire [31:0] dma_dccm_wdata_hi;
	wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_lo;
	wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_hi;
	wire lsu_busm_clken;
	wire lsu_bus_obuf_c1_clken;
	wire lsu_c1_m_clk;
	wire lsu_c1_r_clk;
	wire lsu_c2_m_clk;
	wire lsu_c2_r_clk;
	wire lsu_store_c1_m_clk;
	wire lsu_store_c1_r_clk;
	wire lsu_stbuf_c1_clk;
	wire lsu_bus_ibuf_c1_clk;
	wire lsu_bus_obuf_c1_clk;
	wire lsu_bus_buf_c1_clk;
	wire lsu_busm_clk;
	wire lsu_free_c2_clk;
	wire lsu_raw_fwd_lo_m;
	wire lsu_raw_fwd_hi_m;
	wire lsu_raw_fwd_lo_r;
	wire lsu_raw_fwd_hi_r;
	assign lsu_raw_fwd_lo_m = |stbuf_fwdbyteen_lo_m[pt[1389-:7] - 1:0];
	assign lsu_raw_fwd_hi_m = |stbuf_fwdbyteen_hi_m[pt[1389-:7] - 1:0];
	eb1_lsu_lsc_ctl #(.pt(pt)) lsu_lsc_ctl(
		.rst_l(rst_l),
		.clk_override(clk_override),
		.clk(clk),
		.lsu_c1_m_clk(lsu_c1_m_clk),
		.lsu_c1_r_clk(lsu_c1_r_clk),
		.lsu_c2_m_clk(lsu_c2_m_clk),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.lsu_store_c1_m_clk(lsu_store_c1_m_clk),
		.lsu_ld_data_r(lsu_ld_data_r),
		.lsu_ld_data_corr_r(lsu_ld_data_corr_r),
		.lsu_single_ecc_error_r(lsu_single_ecc_error_r),
		.lsu_double_ecc_error_r(lsu_double_ecc_error_r),
		.lsu_ld_data_m(lsu_ld_data_m),
		.lsu_single_ecc_error_m(lsu_single_ecc_error_m),
		.lsu_double_ecc_error_m(lsu_double_ecc_error_m),
		.flush_m_up(flush_m_up),
		.flush_r(flush_r),
		.ldst_dual_d(ldst_dual_d),
		.ldst_dual_m(ldst_dual_m),
		.ldst_dual_r(ldst_dual_r),
		.exu_lsu_rs1_d(exu_lsu_rs1_d),
		.exu_lsu_rs2_d(exu_lsu_rs2_d),
		.lsu_p(lsu_p),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.dec_lsu_offset_d(dec_lsu_offset_d),
		.picm_mask_data_m(picm_mask_data_m),
		.bus_read_data_m(bus_read_data_m),
		.lsu_result_m(lsu_result_m),
		.lsu_result_corr_r(lsu_result_corr_r),
		.lsu_addr_d(lsu_addr_d),
		.lsu_addr_m(lsu_addr_m),
		.lsu_addr_r(lsu_addr_r),
		.end_addr_d(end_addr_d),
		.end_addr_m(end_addr_m),
		.end_addr_r(end_addr_r),
		.store_data_m(store_data_m),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.lsu_exc_m(lsu_exc_m),
		.is_sideeffects_m(is_sideeffects_m),
		.lsu_commit_r(lsu_commit_r),
		.lsu_single_ecc_error_incr(lsu_single_ecc_error_incr),
		.lsu_error_pkt_r(lsu_error_pkt_r),
		.lsu_fir_addr(lsu_fir_addr),
		.lsu_fir_error(lsu_fir_error),
		.addr_in_dccm_d(addr_in_dccm_d),
		.addr_in_dccm_m(addr_in_dccm_m),
		.addr_in_dccm_r(addr_in_dccm_r),
		.addr_in_pic_d(addr_in_pic_d),
		.addr_in_pic_m(addr_in_pic_m),
		.addr_in_pic_r(addr_in_pic_r),
		.addr_external_m(addr_external_m),
		.dma_dccm_req(dma_dccm_req),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_sz(dma_mem_sz),
		.dma_mem_write(dma_mem_write),
		.dma_mem_wdata(dma_mem_wdata),
		.lsu_pkt_d(lsu_pkt_d),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.scan_mode(scan_mode)
	);
	assign lsu_store_stall_any = (lsu_stbuf_full_any | lsu_bus_buffer_full_any) | ld_single_ecc_error_r_ff;
	assign lsu_load_stall_any = lsu_bus_buffer_full_any | ld_single_ecc_error_r_ff;
	assign lsu_fastint_stall_any = ld_single_ecc_error_r;
	assign dma_mem_tag_d[2:0] = dma_mem_tag[2:0];
	assign ldst_nodma_mtor = ((lsu_pkt_m[0] & ~lsu_pkt_m[4]) & (addr_in_dccm_m | addr_in_pic_m)) & lsu_pkt_m[6];
	assign dccm_ready = ~((dec_lsu_valid_raw_d | ldst_nodma_mtor) | ld_single_ecc_error_r_ff);
	assign dma_dccm_wen = ((dma_dccm_req & dma_mem_write) & addr_in_dccm_d) & dma_mem_sz[1];
	assign dma_pic_wen = (dma_dccm_req & dma_mem_write) & addr_in_pic_d;
	assign {dma_dccm_wdata_hi[31:0], dma_dccm_wdata_lo[31:0]} = dma_mem_wdata[63:0] >> {dma_mem_addr[2:0], 3'b000};
	assign flush_m_up = dec_tlu_flush_lower_r;
	assign flush_r = dec_tlu_i0_kill_writeb_r;
	assign lsu_idle_any = ~((lsu_pkt_m[0] & ~lsu_pkt_m[4]) | (lsu_pkt_r[0] & ~lsu_pkt_r[4])) & lsu_bus_buffer_empty_any;
	assign lsu_active = ((lsu_pkt_m[0] | lsu_pkt_r[0]) | ld_single_ecc_error_r_ff) | ~lsu_bus_buffer_empty_any;
	assign store_stbuf_reqvld_r = (((lsu_pkt_r[0] & lsu_pkt_r[6]) & addr_in_dccm_r) & ~flush_r) & (~lsu_pkt_r[4] | ((lsu_pkt_r[11] | lsu_pkt_r[10]) & ~lsu_double_ecc_error_r));
	assign lsu_cmpen_m = (lsu_pkt_m[0] & (lsu_pkt_m[7] | lsu_pkt_m[6])) & (addr_in_dccm_m | addr_in_pic_m);
	assign lsu_busreq_m = (((lsu_pkt_m[0] & ((lsu_pkt_m[7] | lsu_pkt_m[6]) & addr_external_m)) & ~flush_m_up) & ~lsu_exc_m) & ~lsu_pkt_m[13];
	assign ldst_dual_d = lsu_addr_d[2] != end_addr_d[2];
	assign ldst_dual_m = lsu_addr_m[2] != end_addr_m[2];
	assign ldst_dual_r = lsu_addr_r[2] != end_addr_r[2];
	assign lsu_pmu_misaligned_m = lsu_pkt_m[0] & ((lsu_pkt_m[10] & lsu_addr_m[0]) | (lsu_pkt_m[9] & |lsu_addr_m[1:0]));
	assign lsu_pmu_load_external_m = (lsu_pkt_m[0] & lsu_pkt_m[7]) & addr_external_m;
	assign lsu_pmu_store_external_m = (lsu_pkt_m[0] & lsu_pkt_m[6]) & addr_external_m;
	eb1_lsu_dccm_ctl #(.pt(pt)) dccm_ctl(
		.lsu_addr_d(lsu_addr_d[31:0]),
		.end_addr_d(end_addr_d[pt[1398-:9] - 1:0]),
		.lsu_addr_m(lsu_addr_m[pt[1398-:9] - 1:0]),
		.lsu_addr_r(lsu_addr_r[31:0]),
		.end_addr_m(end_addr_m[pt[1398-:9] - 1:0]),
		.end_addr_r(end_addr_r[pt[1398-:9] - 1:0]),
		.lsu_c2_m_clk(lsu_c2_m_clk),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.lsu_c1_r_clk(lsu_c1_r_clk),
		.lsu_store_c1_r_clk(lsu_store_c1_r_clk),
		.lsu_free_c2_clk(lsu_free_c2_clk),
		.clk_override(clk_override),
		.clk(clk),
		.rst_l(rst_l),
		.lsu_pkt_r(lsu_pkt_r),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_d(lsu_pkt_d),
		.addr_in_dccm_d(addr_in_dccm_d),
		.addr_in_pic_d(addr_in_pic_d),
		.addr_in_pic_m(addr_in_pic_m),
		.addr_in_dccm_m(addr_in_dccm_m),
		.addr_in_dccm_r(addr_in_dccm_r),
		.addr_in_pic_r(addr_in_pic_r),
		.lsu_raw_fwd_lo_r(lsu_raw_fwd_lo_r),
		.lsu_raw_fwd_hi_r(lsu_raw_fwd_hi_r),
		.lsu_commit_r(lsu_commit_r),
		.ldst_dual_m(ldst_dual_m),
		.ldst_dual_r(ldst_dual_r),
		.stbuf_reqvld_any(stbuf_reqvld_any),
		.stbuf_addr_any(stbuf_addr_any),
		.stbuf_data_any(stbuf_data_any),
		.stbuf_ecc_any(stbuf_ecc_any),
		.stbuf_fwddata_hi_m(stbuf_fwddata_hi_m),
		.stbuf_fwddata_lo_m(stbuf_fwddata_lo_m),
		.stbuf_fwdbyteen_hi_m(stbuf_fwdbyteen_hi_m),
		.stbuf_fwdbyteen_lo_m(stbuf_fwdbyteen_lo_m),
		.dccm_rdata_hi_r(dccm_rdata_hi_r),
		.dccm_rdata_lo_r(dccm_rdata_lo_r),
		.dccm_data_ecc_hi_r(dccm_data_ecc_hi_r),
		.dccm_data_ecc_lo_r(dccm_data_ecc_lo_r),
		.lsu_ld_data_r(lsu_ld_data_r),
		.lsu_ld_data_corr_r(lsu_ld_data_corr_r),
		.lsu_double_ecc_error_r(lsu_double_ecc_error_r),
		.single_ecc_error_hi_r(single_ecc_error_hi_r),
		.single_ecc_error_lo_r(single_ecc_error_lo_r),
		.sec_data_hi_r(sec_data_hi_r),
		.sec_data_lo_r(sec_data_lo_r),
		.sec_data_hi_r_ff(sec_data_hi_r_ff),
		.sec_data_lo_r_ff(sec_data_lo_r_ff),
		.sec_data_ecc_hi_r_ff(sec_data_ecc_hi_r_ff),
		.sec_data_ecc_lo_r_ff(sec_data_ecc_lo_r_ff),
		.dccm_rdata_hi_m(dccm_rdata_hi_m),
		.dccm_rdata_lo_m(dccm_rdata_lo_m),
		.dccm_data_ecc_hi_m(dccm_data_ecc_hi_m),
		.dccm_data_ecc_lo_m(dccm_data_ecc_lo_m),
		.lsu_ld_data_m(lsu_ld_data_m),
		.lsu_double_ecc_error_m(lsu_double_ecc_error_m),
		.sec_data_hi_m(sec_data_hi_m),
		.sec_data_lo_m(sec_data_lo_m),
		.store_data_m(store_data_m),
		.dma_dccm_wen(dma_dccm_wen),
		.dma_pic_wen(dma_pic_wen),
		.dma_mem_tag_m(dma_mem_tag_m),
		.dma_mem_addr(dma_mem_addr),
		.dma_mem_wdata(dma_mem_wdata),
		.dma_dccm_wdata_lo(dma_dccm_wdata_lo),
		.dma_dccm_wdata_hi(dma_dccm_wdata_hi),
		.dma_dccm_wdata_ecc_hi(dma_dccm_wdata_ecc_hi),
		.dma_dccm_wdata_ecc_lo(dma_dccm_wdata_ecc_lo),
		.store_data_hi_r(store_data_hi_r),
		.store_data_lo_r(store_data_lo_r),
		.store_datafn_hi_r(store_datafn_hi_r),
		.store_datafn_lo_r(store_datafn_lo_r),
		.store_data_r(store_data_r),
		.ld_single_ecc_error_r(ld_single_ecc_error_r),
		.ld_single_ecc_error_r_ff(ld_single_ecc_error_r_ff),
		.picm_mask_data_m(picm_mask_data_m),
		.lsu_stbuf_commit_any(lsu_stbuf_commit_any),
		.lsu_dccm_rden_m(lsu_dccm_rden_m),
		.lsu_dccm_rden_r(lsu_dccm_rden_r),
		.dccm_dma_rvalid(dccm_dma_rvalid),
		.dccm_dma_ecc_error(dccm_dma_ecc_error),
		.dccm_dma_rtag(dccm_dma_rtag),
		.dccm_dma_rdata(dccm_dma_rdata),
		.dccm_wren(dccm_wren),
		.dccm_rden(dccm_rden),
		.dccm_wr_addr_lo(dccm_wr_addr_lo),
		.dccm_wr_addr_hi(dccm_wr_addr_hi),
		.dccm_rd_addr_lo(dccm_rd_addr_lo),
		.dccm_rd_addr_hi(dccm_rd_addr_hi),
		.dccm_wr_data_lo(dccm_wr_data_lo),
		.dccm_wr_data_hi(dccm_wr_data_hi),
		.dccm_rd_data_lo(dccm_rd_data_lo),
		.dccm_rd_data_hi(dccm_rd_data_hi),
		.picm_wren(picm_wren),
		.picm_rden(picm_rden),
		.picm_mken(picm_mken),
		.picm_rdaddr(picm_rdaddr),
		.picm_wraddr(picm_wraddr),
		.picm_wr_data(picm_wr_data),
		.picm_rd_data(picm_rd_data),
		.scan_mode(scan_mode)
	);
	eb1_lsu_stbuf #(.pt(pt)) stbuf(
		.lsu_addr_d(lsu_addr_d[pt[157-:9] - 1:0]),
		.end_addr_d(end_addr_d[pt[157-:9] - 1:0]),
		.clk(clk),
		.rst_l(rst_l),
		.lsu_stbuf_c1_clk(lsu_stbuf_c1_clk),
		.lsu_free_c2_clk(lsu_free_c2_clk),
		.store_stbuf_reqvld_r(store_stbuf_reqvld_r),
		.lsu_commit_r(lsu_commit_r),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.store_data_hi_r(store_data_hi_r),
		.store_data_lo_r(store_data_lo_r),
		.store_datafn_hi_r(store_datafn_hi_r),
		.store_datafn_lo_r(store_datafn_lo_r),
		.stbuf_reqvld_any(stbuf_reqvld_any),
		.stbuf_reqvld_flushed_any(stbuf_reqvld_flushed_any),
		.stbuf_addr_any(stbuf_addr_any),
		.stbuf_data_any(stbuf_data_any),
		.lsu_stbuf_commit_any(lsu_stbuf_commit_any),
		.lsu_stbuf_full_any(lsu_stbuf_full_any),
		.lsu_stbuf_empty_any(lsu_stbuf_empty_any),
		.ldst_stbuf_reqvld_r(ldst_stbuf_reqvld_r),
		.lsu_addr_m(lsu_addr_m),
		.lsu_addr_r(lsu_addr_r),
		.end_addr_m(end_addr_m),
		.end_addr_r(end_addr_r),
		.ldst_dual_d(ldst_dual_d),
		.ldst_dual_m(ldst_dual_m),
		.ldst_dual_r(ldst_dual_r),
		.addr_in_dccm_m(addr_in_dccm_m),
		.addr_in_dccm_r(addr_in_dccm_r),
		.lsu_cmpen_m(lsu_cmpen_m),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.stbuf_fwddata_hi_m(stbuf_fwddata_hi_m),
		.stbuf_fwddata_lo_m(stbuf_fwddata_lo_m),
		.stbuf_fwdbyteen_hi_m(stbuf_fwdbyteen_hi_m),
		.stbuf_fwdbyteen_lo_m(stbuf_fwdbyteen_lo_m),
		.scan_mode(scan_mode)
	);
	eb1_lsu_ecc #(.pt(pt)) ecc(
		.lsu_addr_r(lsu_addr_r[pt[1398-:9] - 1:0]),
		.end_addr_r(end_addr_r[pt[1398-:9] - 1:0]),
		.lsu_addr_m(lsu_addr_m[pt[1398-:9] - 1:0]),
		.end_addr_m(end_addr_m[pt[1398-:9] - 1:0]),
		.clk(clk),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.clk_override(clk_override),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.stbuf_data_any(stbuf_data_any),
		.dec_tlu_core_ecc_disable(dec_tlu_core_ecc_disable),
		.lsu_dccm_rden_r(lsu_dccm_rden_r),
		.addr_in_dccm_r(addr_in_dccm_r),
		.dccm_rdata_hi_r(dccm_rdata_hi_r),
		.dccm_rdata_lo_r(dccm_rdata_lo_r),
		.dccm_data_ecc_hi_r(dccm_data_ecc_hi_r),
		.dccm_data_ecc_lo_r(dccm_data_ecc_lo_r),
		.sec_data_hi_r(sec_data_hi_r),
		.sec_data_lo_r(sec_data_lo_r),
		.sec_data_hi_r_ff(sec_data_hi_r_ff),
		.sec_data_lo_r_ff(sec_data_lo_r_ff),
		.ld_single_ecc_error_r(ld_single_ecc_error_r),
		.ld_single_ecc_error_r_ff(ld_single_ecc_error_r_ff),
		.lsu_dccm_rden_m(lsu_dccm_rden_m),
		.addr_in_dccm_m(addr_in_dccm_m),
		.dccm_rdata_hi_m(dccm_rdata_hi_m),
		.dccm_rdata_lo_m(dccm_rdata_lo_m),
		.dccm_data_ecc_hi_m(dccm_data_ecc_hi_m),
		.dccm_data_ecc_lo_m(dccm_data_ecc_lo_m),
		.sec_data_hi_m(sec_data_hi_m),
		.sec_data_lo_m(sec_data_lo_m),
		.dma_dccm_wen(dma_dccm_wen),
		.dma_dccm_wdata_lo(dma_dccm_wdata_lo),
		.dma_dccm_wdata_hi(dma_dccm_wdata_hi),
		.dma_dccm_wdata_ecc_hi(dma_dccm_wdata_ecc_hi),
		.dma_dccm_wdata_ecc_lo(dma_dccm_wdata_ecc_lo),
		.stbuf_ecc_any(stbuf_ecc_any),
		.sec_data_ecc_hi_r_ff(sec_data_ecc_hi_r_ff),
		.sec_data_ecc_lo_r_ff(sec_data_ecc_lo_r_ff),
		.single_ecc_error_hi_r(single_ecc_error_hi_r),
		.single_ecc_error_lo_r(single_ecc_error_lo_r),
		.lsu_single_ecc_error_r(lsu_single_ecc_error_r),
		.lsu_double_ecc_error_r(lsu_double_ecc_error_r),
		.lsu_single_ecc_error_m(lsu_single_ecc_error_m),
		.lsu_double_ecc_error_m(lsu_double_ecc_error_m)
	);
	eb1_lsu_trigger #(.pt(pt)) trigger(
		.store_data_m(store_data_m[31:0]),
		.trigger_pkt_any(trigger_pkt_any),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_addr_m(lsu_addr_m),
		.lsu_trigger_match_m(lsu_trigger_match_m)
	);
	eb1_lsu_clkdomain #(.pt(pt)) clkdomain(
		.clk(clk),
		.active_clk(active_clk),
		.rst_l(rst_l),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.clk_override(clk_override),
		.dma_dccm_req(dma_dccm_req),
		.ldst_stbuf_reqvld_r(ldst_stbuf_reqvld_r),
		.stbuf_reqvld_any(stbuf_reqvld_any),
		.stbuf_reqvld_flushed_any(stbuf_reqvld_flushed_any),
		.lsu_busreq_r(lsu_busreq_r),
		.lsu_bus_buffer_pend_any(lsu_bus_buffer_pend_any),
		.lsu_bus_buffer_empty_any(lsu_bus_buffer_empty_any),
		.lsu_stbuf_empty_any(lsu_stbuf_empty_any),
		.lsu_bus_clk_en(lsu_bus_clk_en),
		.lsu_p(lsu_p),
		.lsu_pkt_d(lsu_pkt_d),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.lsu_bus_obuf_c1_clken(lsu_bus_obuf_c1_clken),
		.lsu_busm_clken(lsu_busm_clken),
		.lsu_c1_m_clk(lsu_c1_m_clk),
		.lsu_c1_r_clk(lsu_c1_r_clk),
		.lsu_c2_m_clk(lsu_c2_m_clk),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.lsu_store_c1_m_clk(lsu_store_c1_m_clk),
		.lsu_store_c1_r_clk(lsu_store_c1_r_clk),
		.lsu_stbuf_c1_clk(lsu_stbuf_c1_clk),
		.lsu_bus_obuf_c1_clk(lsu_bus_obuf_c1_clk),
		.lsu_bus_ibuf_c1_clk(lsu_bus_ibuf_c1_clk),
		.lsu_bus_buf_c1_clk(lsu_bus_buf_c1_clk),
		.lsu_busm_clk(lsu_busm_clk),
		.lsu_free_c2_clk(lsu_free_c2_clk),
		.scan_mode(scan_mode)
	);
	eb1_lsu_bus_intf #(.pt(pt)) bus_intf(
		.lsu_addr_m(lsu_addr_m[31:0] & {32 {addr_external_m & lsu_pkt_m[0]}}),
		.lsu_addr_r(lsu_addr_r[31:0] & {32 {lsu_busreq_r}}),
		.end_addr_m(end_addr_m[31:0] & {32 {addr_external_m & lsu_pkt_m[0]}}),
		.end_addr_r(end_addr_r[31:0] & {32 {lsu_busreq_r}}),
		.store_data_r(store_data_r[31:0] & {32 {lsu_busreq_r}}),
		.clk(clk),
		.clk_override(clk_override),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.dec_tlu_external_ldfwd_disable(dec_tlu_external_ldfwd_disable),
		.dec_tlu_wb_coalescing_disable(dec_tlu_wb_coalescing_disable),
		.dec_tlu_sideeffect_posted_disable(dec_tlu_sideeffect_posted_disable),
		.lsu_bus_obuf_c1_clken(lsu_bus_obuf_c1_clken),
		.lsu_busm_clken(lsu_busm_clken),
		.lsu_c1_r_clk(lsu_c1_r_clk),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.lsu_bus_ibuf_c1_clk(lsu_bus_ibuf_c1_clk),
		.lsu_bus_obuf_c1_clk(lsu_bus_obuf_c1_clk),
		.lsu_bus_buf_c1_clk(lsu_bus_buf_c1_clk),
		.lsu_free_c2_clk(lsu_free_c2_clk),
		.active_clk(active_clk),
		.lsu_busm_clk(lsu_busm_clk),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.lsu_busreq_m(lsu_busreq_m),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.lsu_commit_r(lsu_commit_r),
		.is_sideeffects_m(is_sideeffects_m),
		.flush_m_up(flush_m_up),
		.flush_r(flush_r),
		.ldst_dual_d(ldst_dual_d),
		.ldst_dual_m(ldst_dual_m),
		.ldst_dual_r(ldst_dual_r),
		.lsu_busreq_r(lsu_busreq_r),
		.lsu_bus_buffer_pend_any(lsu_bus_buffer_pend_any),
		.lsu_bus_buffer_full_any(lsu_bus_buffer_full_any),
		.lsu_bus_buffer_empty_any(lsu_bus_buffer_empty_any),
		.bus_read_data_m(bus_read_data_m),
		.lsu_imprecise_error_load_any(lsu_imprecise_error_load_any),
		.lsu_imprecise_error_store_any(lsu_imprecise_error_store_any),
		.lsu_imprecise_error_addr_any(lsu_imprecise_error_addr_any),
		.lsu_nonblock_load_valid_m(lsu_nonblock_load_valid_m),
		.lsu_nonblock_load_tag_m(lsu_nonblock_load_tag_m),
		.lsu_nonblock_load_inv_r(lsu_nonblock_load_inv_r),
		.lsu_nonblock_load_inv_tag_r(lsu_nonblock_load_inv_tag_r),
		.lsu_nonblock_load_data_valid(lsu_nonblock_load_data_valid),
		.lsu_nonblock_load_data_error(lsu_nonblock_load_data_error),
		.lsu_nonblock_load_data_tag(lsu_nonblock_load_data_tag),
		.lsu_nonblock_load_data(lsu_nonblock_load_data),
		.lsu_pmu_bus_trxn(lsu_pmu_bus_trxn),
		.lsu_pmu_bus_misaligned(lsu_pmu_bus_misaligned),
		.lsu_pmu_bus_error(lsu_pmu_bus_error),
		.lsu_pmu_bus_busy(lsu_pmu_bus_busy),
		.lsu_axi_awvalid(lsu_axi_awvalid),
		.lsu_axi_awready(lsu_axi_awready),
		.lsu_axi_awid(lsu_axi_awid),
		.lsu_axi_awaddr(lsu_axi_awaddr),
		.lsu_axi_awregion(lsu_axi_awregion),
		.lsu_axi_awlen(lsu_axi_awlen),
		.lsu_axi_awsize(lsu_axi_awsize),
		.lsu_axi_awburst(lsu_axi_awburst),
		.lsu_axi_awlock(lsu_axi_awlock),
		.lsu_axi_awcache(lsu_axi_awcache),
		.lsu_axi_awprot(lsu_axi_awprot),
		.lsu_axi_awqos(lsu_axi_awqos),
		.lsu_axi_wvalid(lsu_axi_wvalid),
		.lsu_axi_wready(lsu_axi_wready),
		.lsu_axi_wdata(lsu_axi_wdata),
		.lsu_axi_wstrb(lsu_axi_wstrb),
		.lsu_axi_wlast(lsu_axi_wlast),
		.lsu_axi_bvalid(lsu_axi_bvalid),
		.lsu_axi_bready(lsu_axi_bready),
		.lsu_axi_bresp(lsu_axi_bresp),
		.lsu_axi_bid(lsu_axi_bid),
		.lsu_axi_arvalid(lsu_axi_arvalid),
		.lsu_axi_arready(lsu_axi_arready),
		.lsu_axi_arid(lsu_axi_arid),
		.lsu_axi_araddr(lsu_axi_araddr),
		.lsu_axi_arregion(lsu_axi_arregion),
		.lsu_axi_arlen(lsu_axi_arlen),
		.lsu_axi_arsize(lsu_axi_arsize),
		.lsu_axi_arburst(lsu_axi_arburst),
		.lsu_axi_arlock(lsu_axi_arlock),
		.lsu_axi_arcache(lsu_axi_arcache),
		.lsu_axi_arprot(lsu_axi_arprot),
		.lsu_axi_arqos(lsu_axi_arqos),
		.lsu_axi_rvalid(lsu_axi_rvalid),
		.lsu_axi_rready(lsu_axi_rready),
		.lsu_axi_rid(lsu_axi_rid),
		.lsu_axi_rdata(lsu_axi_rdata),
		.lsu_axi_rresp(lsu_axi_rresp),
		.lsu_bus_clk_en(lsu_bus_clk_en)
	);
	rvdff #(.WIDTH(3)) dma_mem_tag_mff(
		.rst_l(rst_l),
		.din(dma_mem_tag_d[2:0]),
		.dout(dma_mem_tag_m[2:0]),
		.clk(lsu_c1_m_clk)
	);
	rvdff #(.WIDTH(2)) lsu_raw_fwd_r_ff(
		.rst_l(rst_l),
		.din({lsu_raw_fwd_hi_m, lsu_raw_fwd_lo_m}),
		.dout({lsu_raw_fwd_hi_r, lsu_raw_fwd_lo_r}),
		.clk(lsu_c2_r_clk)
	);
endmodule
module eb1_lsu_addrcheck (
	lsu_c2_m_clk,
	rst_l,
	start_addr_d,
	end_addr_d,
	lsu_pkt_d,
	dec_tlu_mrac_ff,
	rs1_region_d,
	rs1_d,
	is_sideeffects_m,
	addr_in_dccm_d,
	addr_in_pic_d,
	addr_external_d,
	access_fault_d,
	misaligned_fault_d,
	exc_mscause_d,
	fir_dccm_access_error_d,
	fir_nondccm_access_error_d,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire lsu_c2_m_clk;
	input wire rst_l;
	input wire [31:0] start_addr_d;
	input wire [31:0] end_addr_d;
	input wire [13:0] lsu_pkt_d;
	input wire [31:0] dec_tlu_mrac_ff;
	input wire [3:0] rs1_region_d;
	input wire [31:0] rs1_d;
	output wire is_sideeffects_m;
	output wire addr_in_dccm_d;
	output wire addr_in_pic_d;
	output wire addr_external_d;
	output wire access_fault_d;
	output wire misaligned_fault_d;
	output wire [3:0] exc_mscause_d;
	output wire fir_dccm_access_error_d;
	output wire fir_nondccm_access_error_d;
	input wire scan_mode;
	wire non_dccm_access_ok;
	wire is_sideeffects_d;
	wire is_aligned_d;
	wire start_addr_in_dccm_d;
	wire end_addr_in_dccm_d;
	wire start_addr_in_dccm_region_d;
	wire end_addr_in_dccm_region_d;
	wire start_addr_in_pic_d;
	wire end_addr_in_pic_d;
	wire start_addr_in_pic_region_d;
	wire end_addr_in_pic_region_d;
	wire [4:0] csr_idx;
	wire addr_in_iccm;
	wire start_addr_dccm_or_pic;
	wire base_reg_dccm_or_pic;
	wire unmapped_access_fault_d;
	wire mpu_access_fault_d;
	wire picm_access_fault_d;
	wire regpred_access_fault_d;
	wire regcross_misaligned_fault_d;
	wire sideeffect_misaligned_fault_d;
	wire [3:0] access_fault_mscause_d;
	wire [3:0] misaligned_fault_mscause_d;
	generate
		if (pt[1365-:5] == 1) begin : Gen_dccm_enable
			rvrangecheck #(
				.CCM_SADR(pt[1325-:36]),
				.CCM_SIZE(pt[1289-:14])
			) start_addr_dccm_rangecheck(
				.addr(start_addr_d[31:0]),
				.in_range(start_addr_in_dccm_d),
				.in_region(start_addr_in_dccm_region_d)
			);
			rvrangecheck #(
				.CCM_SADR(pt[1325-:36]),
				.CCM_SIZE(pt[1289-:14])
			) end_addr_dccm_rangecheck(
				.addr(end_addr_d[31:0]),
				.in_range(end_addr_in_dccm_d),
				.in_region(end_addr_in_dccm_region_d)
			);
		end
		else begin : Gen_dccm_disable
			assign start_addr_in_dccm_d = 1'b0;
			assign start_addr_in_dccm_region_d = 1'b0;
			assign end_addr_in_dccm_d = 1'b0;
			assign end_addr_in_dccm_region_d = 1'b0;
		end
	endgenerate
	generate
		if (pt[927-:5] == 1) begin : check_iccm
			assign addr_in_iccm = start_addr_d[31:28] == pt[895-:8];
		end
		else assign addr_in_iccm = 1'b0;
	endgenerate
	rvrangecheck #(
		.CCM_SADR(pt[130-:36]),
		.CCM_SIZE(pt[69-:13])
	) start_addr_pic_rangecheck(
		.addr(start_addr_d[31:0]),
		.in_range(start_addr_in_pic_d),
		.in_region(start_addr_in_pic_region_d)
	);
	rvrangecheck #(
		.CCM_SADR(pt[130-:36]),
		.CCM_SIZE(pt[69-:13])
	) end_addr_pic_rangecheck(
		.addr(end_addr_d[31:0]),
		.in_range(end_addr_in_pic_d),
		.in_region(end_addr_in_pic_region_d)
	);
	assign start_addr_dccm_or_pic = start_addr_in_dccm_region_d | start_addr_in_pic_region_d;
	assign base_reg_dccm_or_pic = ((rs1_region_d[3:0] == pt[1333-:8]) & pt[1365-:5]) | (rs1_region_d[3:0] == pt[77-:8]);
	assign addr_in_dccm_d = start_addr_in_dccm_d & end_addr_in_dccm_d;
	assign addr_in_pic_d = start_addr_in_pic_d & end_addr_in_pic_d;
	assign addr_external_d = ~(start_addr_in_dccm_region_d | start_addr_in_pic_region_d);
	assign csr_idx[4:0] = {start_addr_d[31:28], 1'b1};
	assign is_sideeffects_d = ((dec_tlu_mrac_ff[csr_idx] & ~((start_addr_in_dccm_region_d | start_addr_in_pic_region_d) | addr_in_iccm)) & lsu_pkt_d[0]) & (lsu_pkt_d[6] | lsu_pkt_d[7]);
	assign is_aligned_d = ((lsu_pkt_d[9] & (start_addr_d[1:0] == 2'b00)) | (lsu_pkt_d[10] & (start_addr_d[0] == 1'b0))) | lsu_pkt_d[11];
	assign non_dccm_access_ok = ~(|{pt[1733-:5], pt[1728-:5], pt[1723-:5], pt[1718-:5], pt[1713-:5], pt[1708-:5], pt[1703-:5], pt[1698-:5]}) | (((((((((pt[1733-:5] & ((start_addr_d[31:0] | pt[1693-:36]) == (pt[2021-:36] | pt[1693-:36]))) | (pt[1728-:5] & ((start_addr_d[31:0] | pt[1657-:36]) == (pt[1985-:36] | pt[1657-:36])))) | (pt[1723-:5] & ((start_addr_d[31:0] | pt[1621-:36]) == (pt[1949-:36] | pt[1621-:36])))) | (pt[1718-:5] & ((start_addr_d[31:0] | pt[1585-:36]) == (pt[1913-:36] | pt[1585-:36])))) | (pt[1713-:5] & ((start_addr_d[31:0] | pt[1549-:36]) == (pt[1877-:36] | pt[1549-:36])))) | (pt[1708-:5] & ((start_addr_d[31:0] | pt[1513-:36]) == (pt[1841-:36] | pt[1513-:36])))) | (pt[1703-:5] & ((start_addr_d[31:0] | pt[1477-:36]) == (pt[1805-:36] | pt[1477-:36])))) | (pt[1698-:5] & ((start_addr_d[31:0] | pt[1441-:36]) == (pt[1769-:36] | pt[1441-:36])))) & ((((((((pt[1733-:5] & ((end_addr_d[31:0] | pt[1693-:36]) == (pt[2021-:36] | pt[1693-:36]))) | (pt[1728-:5] & ((end_addr_d[31:0] | pt[1657-:36]) == (pt[1985-:36] | pt[1657-:36])))) | (pt[1723-:5] & ((end_addr_d[31:0] | pt[1621-:36]) == (pt[1949-:36] | pt[1621-:36])))) | (pt[1718-:5] & ((end_addr_d[31:0] | pt[1585-:36]) == (pt[1913-:36] | pt[1585-:36])))) | (pt[1713-:5] & ((end_addr_d[31:0] | pt[1549-:36]) == (pt[1877-:36] | pt[1549-:36])))) | (pt[1708-:5] & ((end_addr_d[31:0] | pt[1513-:36]) == (pt[1841-:36] | pt[1513-:36])))) | (pt[1703-:5] & ((end_addr_d[31:0] | pt[1477-:36]) == (pt[1805-:36] | pt[1477-:36])))) | (pt[1698-:5] & ((end_addr_d[31:0] | pt[1441-:36]) == (pt[1769-:36] | pt[1441-:36])))));
	assign regpred_access_fault_d = start_addr_dccm_or_pic ^ base_reg_dccm_or_pic;
	assign picm_access_fault_d = addr_in_pic_d & ((start_addr_d[1:0] != 2'b00) | ~lsu_pkt_d[9]);
	generate
		if (pt[1365-:5] & (pt[1333-:8] == pt[77-:8])) begin
			assign unmapped_access_fault_d = (((start_addr_in_dccm_region_d & ~(start_addr_in_dccm_d | start_addr_in_pic_d)) | (end_addr_in_dccm_region_d & ~(end_addr_in_dccm_d | end_addr_in_pic_d))) | (start_addr_in_dccm_d & end_addr_in_pic_d)) | (start_addr_in_pic_d & end_addr_in_dccm_d);
			assign mpu_access_fault_d = ~start_addr_in_dccm_region_d & ~non_dccm_access_ok;
		end
		else begin
			assign unmapped_access_fault_d = (((start_addr_in_dccm_region_d & ~start_addr_in_dccm_d) | (end_addr_in_dccm_region_d & ~end_addr_in_dccm_d)) | (start_addr_in_pic_region_d & ~start_addr_in_pic_d)) | (end_addr_in_pic_region_d & ~end_addr_in_pic_d);
			assign mpu_access_fault_d = (~start_addr_in_pic_region_d & ~start_addr_in_dccm_region_d) & ~non_dccm_access_ok;
		end
	endgenerate
	assign access_fault_d = ((((unmapped_access_fault_d | mpu_access_fault_d) | picm_access_fault_d) | regpred_access_fault_d) & lsu_pkt_d[0]) & ~lsu_pkt_d[4];
	assign access_fault_mscause_d[3:0] = (unmapped_access_fault_d ? 4'h2 : (mpu_access_fault_d ? 4'h3 : (regpred_access_fault_d ? 4'h5 : (picm_access_fault_d ? 4'h6 : 4'h0))));
	assign regcross_misaligned_fault_d = start_addr_d[31:28] != end_addr_d[31:28];
	assign sideeffect_misaligned_fault_d = is_sideeffects_d & ~is_aligned_d;
	assign misaligned_fault_d = ((regcross_misaligned_fault_d | (sideeffect_misaligned_fault_d & addr_external_d)) & lsu_pkt_d[0]) & ~lsu_pkt_d[4];
	assign misaligned_fault_mscause_d[3:0] = (regcross_misaligned_fault_d ? 4'h2 : (sideeffect_misaligned_fault_d ? 4'h1 : 4'h0));
	assign exc_mscause_d[3:0] = (misaligned_fault_d ? misaligned_fault_mscause_d[3:0] : access_fault_mscause_d[3:0]);
	assign fir_dccm_access_error_d = (((start_addr_in_dccm_region_d & ~start_addr_in_dccm_d) | (end_addr_in_dccm_region_d & ~end_addr_in_dccm_d)) & lsu_pkt_d[0]) & lsu_pkt_d[13];
	assign fir_nondccm_access_error_d = (~(start_addr_in_dccm_region_d & end_addr_in_dccm_region_d) & lsu_pkt_d[0]) & lsu_pkt_d[13];
	rvdff #(.WIDTH(1)) is_sideeffects_mff(
		.din(is_sideeffects_d),
		.dout(is_sideeffects_m),
		.clk(lsu_c2_m_clk),
		.rst_l(rst_l)
	);
endmodule
module eb1_lsu_bus_buffer (
	clk,
	clk_override,
	rst_l,
	scan_mode,
	dec_tlu_external_ldfwd_disable,
	dec_tlu_wb_coalescing_disable,
	dec_tlu_sideeffect_posted_disable,
	dec_tlu_force_halt,
	lsu_bus_obuf_c1_clken,
	lsu_busm_clken,
	lsu_c2_r_clk,
	lsu_bus_ibuf_c1_clk,
	lsu_bus_obuf_c1_clk,
	lsu_bus_buf_c1_clk,
	lsu_free_c2_clk,
	lsu_busm_clk,
	dec_lsu_valid_raw_d,
	lsu_pkt_m,
	lsu_pkt_r,
	lsu_addr_m,
	end_addr_m,
	lsu_addr_r,
	end_addr_r,
	store_data_r,
	no_word_merge_r,
	no_dword_merge_r,
	lsu_busreq_m,
	lsu_busreq_r,
	ld_full_hit_m,
	flush_m_up,
	flush_r,
	lsu_commit_r,
	is_sideeffects_r,
	ldst_dual_d,
	ldst_dual_m,
	ldst_dual_r,
	ldst_byteen_ext_m,
	lsu_bus_buffer_pend_any,
	lsu_bus_buffer_full_any,
	lsu_bus_buffer_empty_any,
	ld_byte_hit_buf_lo,
	ld_byte_hit_buf_hi,
	ld_fwddata_buf_lo,
	ld_fwddata_buf_hi,
	lsu_imprecise_error_load_any,
	lsu_imprecise_error_store_any,
	lsu_imprecise_error_addr_any,
	lsu_nonblock_load_valid_m,
	lsu_nonblock_load_tag_m,
	lsu_nonblock_load_inv_r,
	lsu_nonblock_load_inv_tag_r,
	lsu_nonblock_load_data_valid,
	lsu_nonblock_load_data_error,
	lsu_nonblock_load_data_tag,
	lsu_nonblock_load_data,
	lsu_pmu_bus_trxn,
	lsu_pmu_bus_misaligned,
	lsu_pmu_bus_error,
	lsu_pmu_bus_busy,
	lsu_axi_awvalid,
	lsu_axi_awready,
	lsu_axi_awid,
	lsu_axi_awaddr,
	lsu_axi_awregion,
	lsu_axi_awlen,
	lsu_axi_awsize,
	lsu_axi_awburst,
	lsu_axi_awlock,
	lsu_axi_awcache,
	lsu_axi_awprot,
	lsu_axi_awqos,
	lsu_axi_wvalid,
	lsu_axi_wready,
	lsu_axi_wdata,
	lsu_axi_wstrb,
	lsu_axi_wlast,
	lsu_axi_bvalid,
	lsu_axi_bready,
	lsu_axi_bresp,
	lsu_axi_bid,
	lsu_axi_arvalid,
	lsu_axi_arready,
	lsu_axi_arid,
	lsu_axi_araddr,
	lsu_axi_arregion,
	lsu_axi_arlen,
	lsu_axi_arsize,
	lsu_axi_arburst,
	lsu_axi_arlock,
	lsu_axi_arcache,
	lsu_axi_arprot,
	lsu_axi_arqos,
	lsu_axi_rvalid,
	lsu_axi_rready,
	lsu_axi_rid,
	lsu_axi_rdata,
	lsu_axi_rresp,
	lsu_bus_clk_en,
	lsu_bus_clk_en_q
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire clk_override;
	input wire rst_l;
	input wire scan_mode;
	input wire dec_tlu_external_ldfwd_disable;
	input wire dec_tlu_wb_coalescing_disable;
	input wire dec_tlu_sideeffect_posted_disable;
	input wire dec_tlu_force_halt;
	input wire lsu_bus_obuf_c1_clken;
	input wire lsu_busm_clken;
	input wire lsu_c2_r_clk;
	input wire lsu_bus_ibuf_c1_clk;
	input wire lsu_bus_obuf_c1_clk;
	input wire lsu_bus_buf_c1_clk;
	input wire lsu_free_c2_clk;
	input wire lsu_busm_clk;
	input wire dec_lsu_valid_raw_d;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_r;
	input wire [31:0] lsu_addr_m;
	input wire [31:0] end_addr_m;
	input wire [31:0] lsu_addr_r;
	input wire [31:0] end_addr_r;
	input wire [31:0] store_data_r;
	input wire no_word_merge_r;
	input wire no_dword_merge_r;
	input wire lsu_busreq_m;
	output wire lsu_busreq_r;
	input wire ld_full_hit_m;
	input wire flush_m_up;
	input wire flush_r;
	input wire lsu_commit_r;
	input wire is_sideeffects_r;
	input wire ldst_dual_d;
	input wire ldst_dual_m;
	input wire ldst_dual_r;
	input wire [7:0] ldst_byteen_ext_m;
	output wire lsu_bus_buffer_pend_any;
	output wire lsu_bus_buffer_full_any;
	output wire lsu_bus_buffer_empty_any;
	output wire [3:0] ld_byte_hit_buf_lo;
	output wire [3:0] ld_byte_hit_buf_hi;
	output reg [31:0] ld_fwddata_buf_lo;
	output reg [31:0] ld_fwddata_buf_hi;
	output wire lsu_imprecise_error_load_any;
	output reg lsu_imprecise_error_store_any;
	output wire [31:0] lsu_imprecise_error_addr_any;
	output wire lsu_nonblock_load_valid_m;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	output wire lsu_nonblock_load_inv_r;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	output wire lsu_nonblock_load_data_valid;
	output reg lsu_nonblock_load_data_error;
	output reg [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	output wire [31:0] lsu_nonblock_load_data;
	output wire lsu_pmu_bus_trxn;
	output wire lsu_pmu_bus_misaligned;
	output wire lsu_pmu_bus_error;
	output wire lsu_pmu_bus_busy;
	output wire lsu_axi_awvalid;
	input wire lsu_axi_awready;
	output wire [pt[181-:8] - 1:0] lsu_axi_awid;
	output wire [31:0] lsu_axi_awaddr;
	output wire [3:0] lsu_axi_awregion;
	output wire [7:0] lsu_axi_awlen;
	output wire [2:0] lsu_axi_awsize;
	output wire [1:0] lsu_axi_awburst;
	output wire lsu_axi_awlock;
	output wire [3:0] lsu_axi_awcache;
	output wire [2:0] lsu_axi_awprot;
	output wire [3:0] lsu_axi_awqos;
	output wire lsu_axi_wvalid;
	input wire lsu_axi_wready;
	output wire [63:0] lsu_axi_wdata;
	output wire [7:0] lsu_axi_wstrb;
	output wire lsu_axi_wlast;
	input wire lsu_axi_bvalid;
	output wire lsu_axi_bready;
	input wire [1:0] lsu_axi_bresp;
	input wire [pt[181-:8] - 1:0] lsu_axi_bid;
	output wire lsu_axi_arvalid;
	input wire lsu_axi_arready;
	output wire [pt[181-:8] - 1:0] lsu_axi_arid;
	output wire [31:0] lsu_axi_araddr;
	output wire [3:0] lsu_axi_arregion;
	output wire [7:0] lsu_axi_arlen;
	output wire [2:0] lsu_axi_arsize;
	output wire [1:0] lsu_axi_arburst;
	output wire lsu_axi_arlock;
	output wire [3:0] lsu_axi_arcache;
	output wire [2:0] lsu_axi_arprot;
	output wire [3:0] lsu_axi_arqos;
	input wire lsu_axi_rvalid;
	output wire lsu_axi_rready;
	input wire [pt[181-:8] - 1:0] lsu_axi_rid;
	input wire [63:0] lsu_axi_rdata;
	input wire [1:0] lsu_axi_rresp;
	input wire lsu_bus_clk_en;
	input wire lsu_bus_clk_en_q;
	localparam DEPTH = pt[173-:9];
	localparam DEPTH_LOG2 = pt[164-:7];
	localparam TIMER = 8;
	localparam TIMER_MAX = 7;
	localparam TIMER_LOG2 = 3;
	wire [3:0] ldst_byteen_hi_m;
	wire [3:0] ldst_byteen_lo_m;
	wire [DEPTH - 1:0] ld_addr_hitvec_lo;
	wire [DEPTH - 1:0] ld_addr_hitvec_hi;
	wire [(4 * DEPTH) - 1:0] ld_byte_hitvec_lo;
	wire [(4 * DEPTH) - 1:0] ld_byte_hitvec_hi;
	wire [(4 * DEPTH) - 1:0] ld_byte_hitvecfn_lo;
	wire [(4 * DEPTH) - 1:0] ld_byte_hitvecfn_hi;
	wire ld_addr_ibuf_hit_lo;
	wire ld_addr_ibuf_hit_hi;
	wire [3:0] ld_byte_ibuf_hit_lo;
	wire [3:0] ld_byte_ibuf_hit_hi;
	wire [3:0] ldst_byteen_r;
	wire [3:0] ldst_byteen_hi_r;
	wire [3:0] ldst_byteen_lo_r;
	wire [31:0] store_data_hi_r;
	wire [31:0] store_data_lo_r;
	wire is_aligned_r;
	wire ldst_samedw_r;
	wire lsu_nonblock_load_valid_r;
	reg [31:0] lsu_nonblock_load_data_hi;
	reg [31:0] lsu_nonblock_load_data_lo;
	wire [31:0] lsu_nonblock_data_unalgn;
	wire [1:0] lsu_nonblock_addr_offset;
	wire [1:0] lsu_nonblock_sz;
	wire lsu_nonblock_unsign;
	reg lsu_nonblock_load_data_ready;
	wire [DEPTH - 1:0] CmdPtr0Dec;
	wire [DEPTH - 1:0] CmdPtr1Dec;
	wire [DEPTH - 1:0] RspPtrDec;
	wire [DEPTH_LOG2 - 1:0] CmdPtr0;
	wire [DEPTH_LOG2 - 1:0] CmdPtr1;
	wire [DEPTH_LOG2 - 1:0] RspPtr;
	reg [DEPTH_LOG2 - 1:0] WrPtr0_m;
	wire [DEPTH_LOG2 - 1:0] WrPtr0_r;
	reg [DEPTH_LOG2 - 1:0] WrPtr1_m;
	wire [DEPTH_LOG2 - 1:0] WrPtr1_r;
	reg found_wrptr0;
	reg found_wrptr1;
	wire found_cmdptr0;
	wire found_cmdptr1;
	reg [3:0] buf_numvld_any;
	reg [3:0] buf_numvld_wrcmd_any;
	reg [3:0] buf_numvld_cmd_any;
	reg [3:0] buf_numvld_pend_any;
	reg any_done_wait_state;
	reg bus_sideeffect_pend;
	wire bus_coalescing_disable;
	reg bus_addr_match_pending;
	wire bus_cmd_sent;
	wire bus_cmd_ready;
	wire bus_wcmd_sent;
	wire bus_wdata_sent;
	wire bus_rsp_read;
	wire bus_rsp_write;
	wire [pt[181-:8] - 1:0] bus_rsp_read_tag;
	wire [pt[181-:8] - 1:0] bus_rsp_write_tag;
	wire bus_rsp_read_error;
	wire bus_rsp_write_error;
	wire [63:0] bus_rsp_rdata;
	wire [(DEPTH * 3) - 1:0] buf_state;
	wire [(DEPTH * 2) - 1:0] buf_sz;
	wire [(DEPTH * 32) - 1:0] buf_addr;
	wire [(DEPTH * 4) - 1:0] buf_byteen;
	wire [DEPTH - 1:0] buf_sideeffect;
	wire [DEPTH - 1:0] buf_write;
	wire [DEPTH - 1:0] buf_unsign;
	wire [DEPTH - 1:0] buf_dual;
	wire [DEPTH - 1:0] buf_samedw;
	wire [DEPTH - 1:0] buf_nomerge;
	wire [DEPTH - 1:0] buf_dualhi;
	wire [(DEPTH * DEPTH_LOG2) - 1:0] buf_dualtag;
	wire [DEPTH - 1:0] buf_ldfwd;
	wire [(DEPTH * DEPTH_LOG2) - 1:0] buf_ldfwdtag;
	wire [DEPTH - 1:0] buf_error;
	wire [(DEPTH * 32) - 1:0] buf_data;
	wire [(DEPTH * DEPTH) - 1:0] buf_age;
	wire [(DEPTH * DEPTH) - 1:0] buf_age_younger;
	wire [(DEPTH * DEPTH) - 1:0] buf_rspage;
	wire [(DEPTH * DEPTH) - 1:0] buf_rsp_pickage;
	reg [(DEPTH * 3) - 1:0] buf_nxtstate;
	reg [DEPTH - 1:0] buf_rst;
	reg [DEPTH - 1:0] buf_state_en;
	reg [DEPTH - 1:0] buf_cmd_state_bus_en;
	reg [DEPTH - 1:0] buf_resp_state_bus_en;
	reg [DEPTH - 1:0] buf_state_bus_en;
	wire [DEPTH - 1:0] buf_dual_in;
	wire [DEPTH - 1:0] buf_samedw_in;
	wire [DEPTH - 1:0] buf_nomerge_in;
	wire [DEPTH - 1:0] buf_sideeffect_in;
	wire [DEPTH - 1:0] buf_unsign_in;
	wire [(DEPTH * 2) - 1:0] buf_sz_in;
	wire [DEPTH - 1:0] buf_write_in;
	reg [DEPTH - 1:0] buf_wr_en;
	wire [DEPTH - 1:0] buf_dualhi_in;
	wire [(DEPTH * DEPTH_LOG2) - 1:0] buf_dualtag_in;
	reg [DEPTH - 1:0] buf_ldfwd_en;
	reg [DEPTH - 1:0] buf_ldfwd_in;
	reg [(DEPTH * DEPTH_LOG2) - 1:0] buf_ldfwdtag_in;
	wire [(DEPTH * 4) - 1:0] buf_byteen_in;
	wire [(DEPTH * 32) - 1:0] buf_addr_in;
	reg [(DEPTH * 32) - 1:0] buf_data_in;
	reg [DEPTH - 1:0] buf_error_en;
	reg [DEPTH - 1:0] buf_data_en;
	wire [(DEPTH * DEPTH) - 1:0] buf_age_in;
	wire [(DEPTH * DEPTH) - 1:0] buf_ageQ;
	wire [(DEPTH * DEPTH) - 1:0] buf_rspage_set;
	wire [(DEPTH * DEPTH) - 1:0] buf_rspage_in;
	wire [(DEPTH * DEPTH) - 1:0] buf_rspageQ;
	wire ibuf_valid;
	wire ibuf_dual;
	wire ibuf_samedw;
	wire ibuf_nomerge;
	wire [DEPTH_LOG2 - 1:0] ibuf_tag;
	wire [DEPTH_LOG2 - 1:0] ibuf_dualtag;
	wire ibuf_sideeffect;
	wire ibuf_unsign;
	wire ibuf_write;
	wire [1:0] ibuf_sz;
	wire [3:0] ibuf_byteen;
	wire [31:0] ibuf_addr;
	wire [31:0] ibuf_data;
	wire [2:0] ibuf_timer;
	wire ibuf_byp;
	wire ibuf_wr_en;
	wire ibuf_rst;
	wire ibuf_force_drain;
	wire ibuf_drain_vld;
	wire [DEPTH - 1:0] ibuf_drainvec_vld;
	wire [DEPTH_LOG2 - 1:0] ibuf_tag_in;
	wire [DEPTH_LOG2 - 1:0] ibuf_dualtag_in;
	wire [1:0] ibuf_sz_in;
	wire [31:0] ibuf_addr_in;
	wire [3:0] ibuf_byteen_in;
	wire [31:0] ibuf_data_in;
	wire [2:0] ibuf_timer_in;
	wire [3:0] ibuf_byteen_out;
	wire [31:0] ibuf_data_out;
	wire ibuf_merge_en;
	wire ibuf_merge_in;
	wire obuf_valid;
	wire obuf_write;
	wire obuf_nosend;
	wire obuf_rdrsp_pend;
	wire obuf_sideeffect;
	wire [31:0] obuf_addr;
	wire [63:0] obuf_data;
	wire [1:0] obuf_sz;
	wire [7:0] obuf_byteen;
	wire obuf_merge;
	wire obuf_cmd_done;
	wire obuf_data_done;
	wire [pt[181-:8] - 1:0] obuf_tag0;
	wire [pt[181-:8] - 1:0] obuf_tag1;
	wire [pt[181-:8] - 1:0] obuf_rdrsp_tag;
	wire ibuf_buf_byp;
	wire obuf_force_wr_en;
	wire obuf_wr_wait;
	wire obuf_wr_en;
	wire obuf_wr_enQ;
	wire obuf_rst;
	wire obuf_write_in;
	wire obuf_nosend_in;
	wire obuf_rdrsp_pend_en;
	wire obuf_rdrsp_pend_in;
	wire obuf_sideeffect_in;
	wire obuf_aligned_in;
	wire [31:0] obuf_addr_in;
	wire [63:0] obuf_data_in;
	wire [1:0] obuf_sz_in;
	wire [7:0] obuf_byteen_in;
	wire obuf_merge_in;
	wire obuf_cmd_done_in;
	wire obuf_data_done_in;
	wire [pt[181-:8] - 1:0] obuf_tag0_in;
	wire [pt[181-:8] - 1:0] obuf_tag1_in;
	wire [pt[181-:8] - 1:0] obuf_rdrsp_tag_in;
	wire obuf_merge_en;
	wire [2:0] obuf_wr_timer;
	wire [2:0] obuf_wr_timer_in;
	wire [7:0] obuf_byteen0_in;
	wire [7:0] obuf_byteen1_in;
	wire [63:0] obuf_data0_in;
	wire [63:0] obuf_data1_in;
	wire lsu_axi_awvalid_q;
	wire lsu_axi_awready_q;
	wire lsu_axi_wvalid_q;
	wire lsu_axi_wready_q;
	wire lsu_axi_arvalid_q;
	wire lsu_axi_arready_q;
	wire lsu_axi_bvalid_q;
	wire lsu_axi_bready_q;
	wire lsu_axi_rvalid_q;
	wire lsu_axi_rready_q;
	wire [pt[181-:8] - 1:0] lsu_axi_bid_q;
	wire [pt[181-:8] - 1:0] lsu_axi_rid_q;
	wire [1:0] lsu_axi_bresp_q;
	wire [1:0] lsu_axi_rresp_q;
	reg [pt[181-:8] - 1:0] lsu_imprecise_error_store_tag;
	wire [63:0] lsu_axi_rdata_q;
	function automatic [2:0] f_Enc8to3;
		input reg [7:0] Dec_value;
		reg [2:0] Enc_value;
		begin
			Enc_value[0] = ((Dec_value[1] | Dec_value[3]) | Dec_value[5]) | Dec_value[7];
			Enc_value[1] = ((Dec_value[2] | Dec_value[3]) | Dec_value[6]) | Dec_value[7];
			Enc_value[2] = ((Dec_value[4] | Dec_value[5]) | Dec_value[6]) | Dec_value[7];
			f_Enc8to3 = Enc_value[2:0];
		end
	endfunction
	assign ldst_byteen_hi_m[3:0] = ldst_byteen_ext_m[7:4];
	assign ldst_byteen_lo_m[3:0] = ldst_byteen_ext_m[3:0];
	localparam [2:0] IDLE = 3'b000;
	generate
		genvar i;
		for (i = 0; i < DEPTH; i = i + 1) begin
			assign ld_addr_hitvec_lo[i] = (((lsu_addr_m[31:2] == buf_addr[(i * 32) + 31-:30]) & buf_write[i]) & (buf_state[i * 3+:3] != IDLE)) & lsu_busreq_m;
			assign ld_addr_hitvec_hi[i] = (((end_addr_m[31:2] == buf_addr[(i * 32) + 31-:30]) & buf_write[i]) & (buf_state[i * 3+:3] != IDLE)) & lsu_busreq_m;
		end
	endgenerate
	generate
		genvar j;
		for (j = 0; j < 4; j = j + 1) begin
			assign ld_byte_hit_buf_lo[j] = |ld_byte_hitvecfn_lo[j * DEPTH+:DEPTH] | ld_byte_ibuf_hit_lo[j];
			assign ld_byte_hit_buf_hi[j] = |ld_byte_hitvecfn_hi[j * DEPTH+:DEPTH] | ld_byte_ibuf_hit_hi[j];
			for (i = 0; i < DEPTH; i = i + 1) begin
				assign ld_byte_hitvec_lo[(j * DEPTH) + i] = (ld_addr_hitvec_lo[i] & buf_byteen[(i * 4) + j]) & ldst_byteen_lo_m[j];
				assign ld_byte_hitvec_hi[(j * DEPTH) + i] = (ld_addr_hitvec_hi[i] & buf_byteen[(i * 4) + j]) & ldst_byteen_hi_m[j];
				assign ld_byte_hitvecfn_lo[(j * DEPTH) + i] = (ld_byte_hitvec_lo[(j * DEPTH) + i] & ~(|(ld_byte_hitvec_lo[j * DEPTH+:DEPTH] & buf_age_younger[i * DEPTH+:DEPTH]))) & ~ld_byte_ibuf_hit_lo[j];
				assign ld_byte_hitvecfn_hi[(j * DEPTH) + i] = (ld_byte_hitvec_hi[(j * DEPTH) + i] & ~(|(ld_byte_hitvec_hi[j * DEPTH+:DEPTH] & buf_age_younger[i * DEPTH+:DEPTH]))) & ~ld_byte_ibuf_hit_hi[j];
			end
		end
	endgenerate
	assign ld_addr_ibuf_hit_lo = (((lsu_addr_m[31:2] == ibuf_addr[31:2]) & ibuf_write) & ibuf_valid) & lsu_busreq_m;
	assign ld_addr_ibuf_hit_hi = (((end_addr_m[31:2] == ibuf_addr[31:2]) & ibuf_write) & ibuf_valid) & lsu_busreq_m;
	generate
		for (i = 0; i < 4; i = i + 1) begin
			assign ld_byte_ibuf_hit_lo[i] = (ld_addr_ibuf_hit_lo & ibuf_byteen[i]) & ldst_byteen_lo_m[i];
			assign ld_byte_ibuf_hit_hi[i] = (ld_addr_ibuf_hit_hi & ibuf_byteen[i]) & ldst_byteen_hi_m[i];
		end
	endgenerate
	always @(*) begin
		ld_fwddata_buf_lo[31:0] = {{8 {ld_byte_ibuf_hit_lo[3]}}, {8 {ld_byte_ibuf_hit_lo[2]}}, {8 {ld_byte_ibuf_hit_lo[1]}}, {8 {ld_byte_ibuf_hit_lo[0]}}} & ibuf_data[31:0];
		ld_fwddata_buf_hi[31:0] = {{8 {ld_byte_ibuf_hit_hi[3]}}, {8 {ld_byte_ibuf_hit_hi[2]}}, {8 {ld_byte_ibuf_hit_hi[1]}}, {8 {ld_byte_ibuf_hit_hi[0]}}} & ibuf_data[31:0];
		begin : sv2v_autoblock_50
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					ld_fwddata_buf_lo[7:0] = ld_fwddata_buf_lo[7:0] | ({8 {ld_byte_hitvecfn_lo[i]}} & buf_data[(i * 32) + 7-:8]);
					ld_fwddata_buf_lo[15:8] = ld_fwddata_buf_lo[15:8] | ({8 {ld_byte_hitvecfn_lo[DEPTH + i]}} & buf_data[(i * 32) + 15-:8]);
					ld_fwddata_buf_lo[23:16] = ld_fwddata_buf_lo[23:16] | ({8 {ld_byte_hitvecfn_lo[(2 * DEPTH) + i]}} & buf_data[(i * 32) + 23-:8]);
					ld_fwddata_buf_lo[31:24] = ld_fwddata_buf_lo[31:24] | ({8 {ld_byte_hitvecfn_lo[(3 * DEPTH) + i]}} & buf_data[(i * 32) + 31-:8]);
					ld_fwddata_buf_hi[7:0] = ld_fwddata_buf_hi[7:0] | ({8 {ld_byte_hitvecfn_hi[i]}} & buf_data[(i * 32) + 7-:8]);
					ld_fwddata_buf_hi[15:8] = ld_fwddata_buf_hi[15:8] | ({8 {ld_byte_hitvecfn_hi[DEPTH + i]}} & buf_data[(i * 32) + 15-:8]);
					ld_fwddata_buf_hi[23:16] = ld_fwddata_buf_hi[23:16] | ({8 {ld_byte_hitvecfn_hi[(2 * DEPTH) + i]}} & buf_data[(i * 32) + 23-:8]);
					ld_fwddata_buf_hi[31:24] = ld_fwddata_buf_hi[31:24] | ({8 {ld_byte_hitvecfn_hi[(3 * DEPTH) + i]}} & buf_data[(i * 32) + 31-:8]);
				end
		end
	end
	assign bus_coalescing_disable = dec_tlu_wb_coalescing_disable | pt[2038];
	assign ldst_byteen_r[3:0] = (({4 {lsu_pkt_r[11]}} & 4'b0001) | ({4 {lsu_pkt_r[10]}} & 4'b0011)) | ({4 {lsu_pkt_r[9]}} & 4'b1111);
	assign {ldst_byteen_hi_r[3:0], ldst_byteen_lo_r[3:0]} = {4'b0000, ldst_byteen_r[3:0]} << lsu_addr_r[1:0];
	assign {store_data_hi_r[31:0], store_data_lo_r[31:0]} = {32'b00000000000000000000000000000000, store_data_r[31:0]} << (8 * lsu_addr_r[1:0]);
	assign ldst_samedw_r = lsu_addr_r[3] == end_addr_r[3];
	assign is_aligned_r = ((lsu_pkt_r[9] & (lsu_addr_r[1:0] == 2'b00)) | (lsu_pkt_r[10] & (lsu_addr_r[0] == 1'b0))) | lsu_pkt_r[11];
	assign ibuf_byp = (lsu_busreq_r & (lsu_pkt_r[7] | no_word_merge_r)) & ~ibuf_valid;
	assign ibuf_wr_en = (lsu_busreq_r & lsu_commit_r) & ~ibuf_byp;
	assign ibuf_rst = (ibuf_drain_vld & ~ibuf_wr_en) | dec_tlu_force_halt;
	assign ibuf_force_drain = ((lsu_busreq_m & ~lsu_busreq_r) & ibuf_valid) & (lsu_pkt_m[7] | (ibuf_addr[31:2] != lsu_addr_m[31:2]));
	assign ibuf_drain_vld = ibuf_valid & (((((((ibuf_wr_en | (ibuf_timer == TIMER_MAX)) & ~(ibuf_merge_en & ibuf_merge_in)) | ibuf_byp) | ibuf_force_drain) | ibuf_sideeffect) | ~ibuf_write) | bus_coalescing_disable);
	assign ibuf_tag_in[DEPTH_LOG2 - 1:0] = (ibuf_merge_en & ibuf_merge_in ? ibuf_tag[DEPTH_LOG2 - 1:0] : (ldst_dual_r ? WrPtr1_r : WrPtr0_r));
	assign ibuf_dualtag_in[DEPTH_LOG2 - 1:0] = WrPtr0_r;
	assign ibuf_sz_in[1:0] = {lsu_pkt_r[9], lsu_pkt_r[10]};
	assign ibuf_addr_in[31:0] = (ldst_dual_r ? end_addr_r[31:0] : lsu_addr_r[31:0]);
	assign ibuf_byteen_in[3:0] = (ibuf_merge_en & ibuf_merge_in ? ibuf_byteen[3:0] | ldst_byteen_lo_r[3:0] : (ldst_dual_r ? ldst_byteen_hi_r[3:0] : ldst_byteen_lo_r[3:0]));
	generate
		for (i = 0; i < 4; i = i + 1) assign ibuf_data_in[(8 * i) + 7:8 * i] = (ibuf_merge_en & ibuf_merge_in ? (ldst_byteen_lo_r[i] ? store_data_lo_r[(8 * i) + 7:8 * i] : ibuf_data[(8 * i) + 7:8 * i]) : (ldst_dual_r ? store_data_hi_r[(8 * i) + 7:8 * i] : store_data_lo_r[(8 * i) + 7:8 * i]));
	endgenerate
	assign ibuf_timer_in = (ibuf_wr_en ? {3 {1'sb0}} : (ibuf_timer < TIMER_MAX ? ibuf_timer + 1'b1 : ibuf_timer));
	assign ibuf_merge_en = ((((((lsu_busreq_r & lsu_commit_r) & lsu_pkt_r[6]) & ibuf_valid) & ibuf_write) & (lsu_addr_r[31:2] == ibuf_addr[31:2])) & ~is_sideeffects_r) & ~bus_coalescing_disable;
	assign ibuf_merge_in = ~ldst_dual_r;
	generate
		for (i = 0; i < 4; i = i + 1) begin
			assign ibuf_byteen_out[i] = (ibuf_merge_en & ~ibuf_merge_in ? ibuf_byteen[i] | ldst_byteen_lo_r[i] : ibuf_byteen[i]);
			assign ibuf_data_out[(8 * i) + 7:8 * i] = (ibuf_merge_en & ~ibuf_merge_in ? (ldst_byteen_lo_r[i] ? store_data_lo_r[(8 * i) + 7:8 * i] : ibuf_data[(8 * i) + 7:8 * i]) : ibuf_data[(8 * i) + 7:8 * i]);
		end
	endgenerate
	rvdffsc #(.WIDTH(1)) ibuf_valid_ff(
		.din(1'b1),
		.dout(ibuf_valid),
		.en(ibuf_wr_en),
		.clear(ibuf_rst),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(DEPTH_LOG2)) ibuf_tagff(
		.din(ibuf_tag_in),
		.dout(ibuf_tag),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(DEPTH_LOG2)) ibuf_dualtagff(
		.din(ibuf_dualtag_in),
		.dout(ibuf_dualtag),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_dualff(
		.din(ldst_dual_r),
		.dout(ibuf_dual),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_samedwff(
		.din(ldst_samedw_r),
		.dout(ibuf_samedw),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_nomergeff(
		.din(no_dword_merge_r),
		.dout(ibuf_nomerge),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_sideeffectff(
		.din(is_sideeffects_r),
		.dout(ibuf_sideeffect),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_unsignff(
		.din(lsu_pkt_r[5]),
		.dout(ibuf_unsign),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) ibuf_writeff(
		.din(lsu_pkt_r[6]),
		.dout(ibuf_write),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(2)) ibuf_szff(
		.din(ibuf_sz_in[1:0]),
		.dout(ibuf_sz),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) ibuf_addrff(
		.din(ibuf_addr_in[31:0]),
		.dout(ibuf_addr),
		.en(ibuf_wr_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffs #(.WIDTH(4)) ibuf_byteenff(
		.din(ibuf_byteen_in[3:0]),
		.dout(ibuf_byteen),
		.en(ibuf_wr_en),
		.clk(lsu_bus_ibuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) ibuf_dataff(
		.din(ibuf_data_in[31:0]),
		.dout(ibuf_data),
		.en(ibuf_wr_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdff #(.WIDTH(TIMER_LOG2)) ibuf_timerff(
		.din(ibuf_timer_in),
		.dout(ibuf_timer),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	assign obuf_wr_wait = ((((((buf_numvld_wrcmd_any[3:0] == 4'b0001) & (buf_numvld_cmd_any[3:0] == 4'b0001)) & (obuf_wr_timer != TIMER_MAX)) & ~bus_coalescing_disable) & ~buf_nomerge[CmdPtr0]) & ~buf_sideeffect[CmdPtr0]) & ~obuf_force_wr_en;
	assign obuf_wr_timer_in = (obuf_wr_en ? 3'b000 : ((buf_numvld_cmd_any > 4'b0000) & (obuf_wr_timer < TIMER_MAX) ? obuf_wr_timer + 1'b1 : obuf_wr_timer));
	assign obuf_force_wr_en = (((lsu_busreq_m & ~lsu_busreq_r) & ~ibuf_valid) & (buf_numvld_cmd_any[3:0] == 4'b0001)) & (lsu_addr_m[31:2] != buf_addr[(CmdPtr0 * 32) + 31-:30]);
	assign ibuf_buf_byp = (ibuf_byp & (buf_numvld_pend_any[3:0] == 4'b0000)) & (~lsu_pkt_r[6] | no_dword_merge_r);
	localparam [2:0] CMD = 3'b010;
	assign obuf_wr_en = ((((((ibuf_buf_byp & lsu_commit_r) & ~(is_sideeffects_r & bus_sideeffect_pend)) | (((((buf_state[CmdPtr0 * 3+:3] == CMD) & found_cmdptr0) & ~buf_cmd_state_bus_en[CmdPtr0]) & ~(buf_sideeffect[CmdPtr0] & bus_sideeffect_pend)) & (((~((buf_dual[CmdPtr0] & buf_samedw[CmdPtr0]) & ~buf_write[CmdPtr0]) | found_cmdptr1) | buf_nomerge[CmdPtr0]) | obuf_force_wr_en))) & ((bus_cmd_ready | ~obuf_valid) | obuf_nosend)) & ~obuf_wr_wait) & ~bus_addr_match_pending) & lsu_bus_clk_en;
	assign obuf_rst = (((bus_cmd_sent | (obuf_valid & obuf_nosend)) & ~obuf_wr_en) & lsu_bus_clk_en) | dec_tlu_force_halt;
	assign obuf_write_in = (ibuf_buf_byp ? lsu_pkt_r[6] : buf_write[CmdPtr0]);
	assign obuf_sideeffect_in = (ibuf_buf_byp ? is_sideeffects_r : buf_sideeffect[CmdPtr0]);
	assign obuf_addr_in[31:0] = (ibuf_buf_byp ? lsu_addr_r[31:0] : buf_addr[CmdPtr0 * 32+:32]);
	assign obuf_sz_in[1:0] = (ibuf_buf_byp ? {lsu_pkt_r[9], lsu_pkt_r[10]} : buf_sz[CmdPtr0 * 2+:2]);
	assign obuf_merge_in = obuf_merge_en;
	function automatic [pt[181-:8] - 1:0] sv2v_cast_72B45;
		input reg [pt[181-:8] - 1:0] inp;
		sv2v_cast_72B45 = inp;
	endfunction
	assign obuf_tag0_in[pt[181-:8] - 1:0] = (ibuf_buf_byp ? sv2v_cast_72B45(WrPtr0_r) : sv2v_cast_72B45(CmdPtr0));
	assign obuf_tag1_in[pt[181-:8] - 1:0] = (ibuf_buf_byp ? sv2v_cast_72B45(WrPtr1_r) : sv2v_cast_72B45(CmdPtr1));
	assign obuf_cmd_done_in = ~(obuf_wr_en | obuf_rst) & (obuf_cmd_done | bus_wcmd_sent);
	assign obuf_data_done_in = ~(obuf_wr_en | obuf_rst) & (obuf_data_done | bus_wdata_sent);
	assign obuf_aligned_in = (ibuf_buf_byp ? is_aligned_r : ((obuf_sz_in[1:0] == 2'b00) | (obuf_sz_in[0] & ~obuf_addr_in[0])) | (obuf_sz_in[1] & ~(|obuf_addr_in[1:0])));
	assign obuf_rdrsp_pend_in = (((~(obuf_wr_en & ~obuf_nosend_in) & obuf_rdrsp_pend) & ~(bus_rsp_read & (bus_rsp_read_tag == obuf_rdrsp_tag))) | (bus_cmd_sent & ~obuf_write)) & ~dec_tlu_force_halt;
	assign obuf_rdrsp_pend_en = lsu_bus_clk_en | dec_tlu_force_halt;
	assign obuf_rdrsp_tag_in[pt[181-:8] - 1:0] = (bus_cmd_sent & ~obuf_write ? obuf_tag0[pt[181-:8] - 1:0] : obuf_rdrsp_tag[pt[181-:8] - 1:0]);
	assign obuf_nosend_in = ((((((obuf_addr_in[31:3] == obuf_addr[31:3]) & obuf_aligned_in) & ~obuf_sideeffect) & ~obuf_write) & ~obuf_write_in) & ~dec_tlu_external_ldfwd_disable) & ((obuf_valid & ~obuf_nosend) | (obuf_rdrsp_pend & ~(bus_rsp_read & (bus_rsp_read_tag == obuf_rdrsp_tag))));
	assign obuf_byteen0_in[7:0] = (ibuf_buf_byp ? (lsu_addr_r[2] ? {ldst_byteen_lo_r[3:0], 4'b0000} : {4'b0000, ldst_byteen_lo_r[3:0]}) : (buf_addr[(CmdPtr0 * 32) + 2] ? {buf_byteen[CmdPtr0 * 4+:4], 4'b0000} : {4'b0000, buf_byteen[CmdPtr0 * 4+:4]}));
	assign obuf_byteen1_in[7:0] = (ibuf_buf_byp ? (end_addr_r[2] ? {ldst_byteen_hi_r[3:0], 4'b0000} : {4'b0000, ldst_byteen_hi_r[3:0]}) : (buf_addr[(CmdPtr1 * 32) + 2] ? {buf_byteen[CmdPtr1 * 4+:4], 4'b0000} : {4'b0000, buf_byteen[CmdPtr1 * 4+:4]}));
	assign obuf_data0_in[63:0] = (ibuf_buf_byp ? (lsu_addr_r[2] ? {store_data_lo_r[31:0], 32'b00000000000000000000000000000000} : {32'b00000000000000000000000000000000, store_data_lo_r[31:0]}) : (buf_addr[(CmdPtr0 * 32) + 2] ? {buf_data[CmdPtr0 * 32+:32], 32'b00000000000000000000000000000000} : {32'b00000000000000000000000000000000, buf_data[CmdPtr0 * 32+:32]}));
	assign obuf_data1_in[63:0] = (ibuf_buf_byp ? (end_addr_r[2] ? {store_data_hi_r[31:0], 32'b00000000000000000000000000000000} : {32'b00000000000000000000000000000000, store_data_hi_r[31:0]}) : (buf_addr[(CmdPtr1 * 32) + 2] ? {buf_data[CmdPtr1 * 32+:32], 32'b00000000000000000000000000000000} : {32'b00000000000000000000000000000000, buf_data[CmdPtr1 * 32+:32]}));
	generate
		for (i = 0; i < 8; i = i + 1) begin
			assign obuf_byteen_in[i] = obuf_byteen0_in[i] | (obuf_merge_en & obuf_byteen1_in[i]);
			assign obuf_data_in[(8 * i) + 7:8 * i] = (obuf_merge_en & obuf_byteen1_in[i] ? obuf_data1_in[(8 * i) + 7:8 * i] : obuf_data0_in[(8 * i) + 7:8 * i]);
		end
	endgenerate
	assign obuf_merge_en = ((((((((CmdPtr0 != CmdPtr1) & found_cmdptr0) & found_cmdptr1) & (buf_state[CmdPtr0 * 3+:3] == CMD)) & (buf_state[CmdPtr1 * 3+:3] == CMD)) & ~buf_cmd_state_bus_en[CmdPtr0]) & ~buf_sideeffect[CmdPtr0]) & (((~buf_write[CmdPtr0] & buf_dual[CmdPtr0]) & ~buf_dualhi[CmdPtr0]) & buf_samedw[CmdPtr0])) | ((ibuf_buf_byp & ldst_samedw_r) & ldst_dual_r);
	rvdff_fpga #(.WIDTH(1)) obuf_wren_ff(
		.din(obuf_wr_en),
		.dout(obuf_wr_enQ),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffsc #(.WIDTH(1)) obuf_valid_ff(
		.din(1'b1),
		.dout(obuf_valid),
		.en(obuf_wr_en),
		.clear(obuf_rst),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) obuf_nosend_ff(
		.din(obuf_nosend_in),
		.dout(obuf_nosend),
		.en(obuf_wr_en),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(1)) obuf_rdrsp_pend_ff(
		.din(obuf_rdrsp_pend_in),
		.dout(obuf_rdrsp_pend),
		.en(obuf_rdrsp_pend_en),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) obuf_cmd_done_ff(
		.din(obuf_cmd_done_in),
		.dout(obuf_cmd_done),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) obuf_data_done_ff(
		.din(obuf_data_done_in),
		.dout(obuf_data_done),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(pt[181-:8])) obuf_rdrsp_tagff(
		.din(obuf_rdrsp_tag_in),
		.dout(obuf_rdrsp_tag),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(pt[181-:8])) obuf_tag0ff(
		.din(obuf_tag0_in),
		.dout(obuf_tag0),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(pt[181-:8])) obuf_tag1ff(
		.din(obuf_tag1_in),
		.dout(obuf_tag1),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) obuf_mergeff(
		.din(obuf_merge_in),
		.dout(obuf_merge),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) obuf_writeff(
		.din(obuf_write_in),
		.dout(obuf_write),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(1)) obuf_sideeffectff(
		.din(obuf_sideeffect_in),
		.dout(obuf_sideeffect),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(2)) obuf_szff(
		.din(obuf_sz_in[1:0]),
		.dout(obuf_sz),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffs_fpga #(.WIDTH(8)) obuf_byteenff(
		.din(obuf_byteen_in[7:0]),
		.dout(obuf_byteen),
		.en(obuf_wr_en),
		.clk(lsu_bus_obuf_c1_clk),
		.clken(lsu_bus_obuf_c1_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) obuf_addrff(
		.din(obuf_addr_in[31:0]),
		.dout(obuf_addr),
		.en(obuf_wr_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffe #(.WIDTH(64)) obuf_dataff(
		.din(obuf_data_in[63:0]),
		.dout(obuf_data),
		.en(obuf_wr_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdff_fpga #(.WIDTH(TIMER_LOG2)) obuf_timerff(
		.din(obuf_wr_timer_in),
		.dout(obuf_wr_timer),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	function automatic signed [DEPTH_LOG2 - 1:0] sv2v_cast_63A9F_signed;
		input reg signed [DEPTH_LOG2 - 1:0] inp;
		sv2v_cast_63A9F_signed = inp;
	endfunction
	always @(*) begin
		WrPtr0_m[DEPTH_LOG2 - 1:0] = {DEPTH_LOG2 {1'sb0}};
		WrPtr1_m[DEPTH_LOG2 - 1:0] = {DEPTH_LOG2 {1'sb0}};
		found_wrptr0 = 1'b0;
		found_wrptr1 = 1'b0;
		begin : sv2v_autoblock_51
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				if (~found_wrptr0) begin
					WrPtr0_m[DEPTH_LOG2 - 1:0] = sv2v_cast_63A9F_signed(i);
					found_wrptr0 = (buf_state[i * 3+:3] == IDLE) & ~((ibuf_valid & (ibuf_tag == i)) | (lsu_busreq_r & ((WrPtr0_r == i) | (ldst_dual_r & (WrPtr1_r == i)))));
				end
		end
		begin : sv2v_autoblock_52
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				if (~found_wrptr1) begin
					WrPtr1_m[DEPTH_LOG2 - 1:0] = sv2v_cast_63A9F_signed(i);
					found_wrptr1 = (buf_state[i * 3+:3] == IDLE) & ~(((ibuf_valid & (ibuf_tag == i)) | (lsu_busreq_m & (WrPtr0_m == i))) | (lsu_busreq_r & ((WrPtr0_r == i) | (ldst_dual_r & (WrPtr1_r == i)))));
				end
		end
	end
	localparam [2:0] DONE_WAIT = 3'b101;
	generate
		for (i = 0; i < DEPTH; i = i + 1) begin
			assign CmdPtr0Dec[i] = (~(|buf_age[i * DEPTH+:DEPTH]) & (buf_state[i * 3+:3] == CMD)) & ~buf_cmd_state_bus_en[i];
			assign CmdPtr1Dec[i] = ((~(|(buf_age[i * DEPTH+:DEPTH] & ~CmdPtr0Dec)) & ~CmdPtr0Dec[i]) & (buf_state[i * 3+:3] == CMD)) & ~buf_cmd_state_bus_en[i];
			assign RspPtrDec[i] = ~(|buf_rsp_pickage[i * DEPTH+:DEPTH]) & (buf_state[i * 3+:3] == DONE_WAIT);
		end
	endgenerate
	assign found_cmdptr0 = |CmdPtr0Dec;
	assign found_cmdptr1 = |CmdPtr1Dec;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	assign CmdPtr0 = f_Enc8to3(sv2v_cast_8(CmdPtr0Dec[DEPTH - 1:0]));
	assign CmdPtr1 = f_Enc8to3(sv2v_cast_8(CmdPtr1Dec[DEPTH - 1:0]));
	assign RspPtr = f_Enc8to3(sv2v_cast_8(RspPtrDec[DEPTH - 1:0]));
	localparam [2:0] WAIT = 3'b001;
	generate
		for (i = 0; i < DEPTH; i = i + 1) begin : GenAgeVec
			for (j = 0; j < DEPTH; j = j + 1) begin
				assign buf_age_in[(i * DEPTH) + j] = (((buf_state[i * 3+:3] == IDLE) & buf_state_en[i]) & ((((buf_state[j * 3+:3] == WAIT) | ((buf_state[j * 3+:3] == CMD) & ~buf_cmd_state_bus_en[j])) | ((((ibuf_drain_vld & lsu_busreq_r) & (ibuf_byp | ldst_dual_r)) & (i == WrPtr0_r)) & (j == ibuf_tag))) | ((((ibuf_byp & lsu_busreq_r) & ldst_dual_r) & (i == WrPtr1_r)) & (j == WrPtr0_r)))) | buf_age[(i * DEPTH) + j];
				assign buf_age[(i * DEPTH) + j] = (buf_ageQ[(i * DEPTH) + j] & ~((buf_state[j * 3+:3] == CMD) & buf_cmd_state_bus_en[j])) & ~dec_tlu_force_halt;
				assign buf_age_younger[(i * DEPTH) + j] = (i == j ? 1'b0 : ~buf_age[(i * DEPTH) + j] & (buf_state[j * 3+:3] != IDLE));
			end
		end
	endgenerate
	localparam [2:0] DONE = 3'b110;
	generate
		for (i = 0; i < DEPTH; i = i + 1) begin : GenRspAgeVec
			for (j = 0; j < DEPTH; j = j + 1) begin
				function automatic signed [DEPTH_LOG2 - 1:0] sv2v_cast_63A9F_signed;
					input reg signed [DEPTH_LOG2 - 1:0] inp;
					sv2v_cast_63A9F_signed = inp;
				endfunction
				assign buf_rspage_set[(i * DEPTH) + j] = ((buf_state[i * 3+:3] == IDLE) & buf_state_en[i]) & ((~((buf_state[j * 3+:3] == IDLE) | (buf_state[j * 3+:3] == DONE)) | ((((ibuf_drain_vld & lsu_busreq_r) & (ibuf_byp | ldst_dual_r)) & (sv2v_cast_63A9F_signed(i) == WrPtr0_r)) & (sv2v_cast_63A9F_signed(j) == ibuf_tag))) | ((((ibuf_byp & lsu_busreq_r) & ldst_dual_r) & (sv2v_cast_63A9F_signed(i) == WrPtr1_r)) & (sv2v_cast_63A9F_signed(j) == WrPtr0_r)));
				assign buf_rspage_in[(i * DEPTH) + j] = buf_rspage_set[(i * DEPTH) + j] | buf_rspage[(i * DEPTH) + j];
				assign buf_rspage[(i * DEPTH) + j] = (buf_rspageQ[(i * DEPTH) + j] & ~((buf_state[j * 3+:3] == DONE) | (buf_state[j * 3+:3] == IDLE))) & ~dec_tlu_force_halt;
				assign buf_rsp_pickage[(i * DEPTH) + j] = buf_rspageQ[(i * DEPTH) + j] & (buf_state[j * 3+:3] == DONE_WAIT);
			end
		end
	endgenerate
	localparam [2:0] DONE_PARTIAL = 3'b100;
	localparam [2:0] RESP = 3'b011;
	generate
		for (i = 0; i < DEPTH; i = i + 1) begin
			assign ibuf_drainvec_vld[i] = ibuf_drain_vld & (i == ibuf_tag);
			assign buf_byteen_in[i * 4+:4] = (ibuf_drainvec_vld[i] ? ibuf_byteen_out[3:0] : ((ibuf_byp & ldst_dual_r) & (i == WrPtr1_r) ? ldst_byteen_hi_r[3:0] : ldst_byteen_lo_r[3:0]));
			assign buf_addr_in[i * 32+:32] = (ibuf_drainvec_vld[i] ? ibuf_addr[31:0] : ((ibuf_byp & ldst_dual_r) & (i == WrPtr1_r) ? end_addr_r[31:0] : lsu_addr_r[31:0]));
			assign buf_dual_in[i] = (ibuf_drainvec_vld[i] ? ibuf_dual : ldst_dual_r);
			assign buf_samedw_in[i] = (ibuf_drainvec_vld[i] ? ibuf_samedw : ldst_samedw_r);
			assign buf_nomerge_in[i] = (ibuf_drainvec_vld[i] ? ibuf_nomerge | ibuf_force_drain : no_dword_merge_r);
			assign buf_dualhi_in[i] = (ibuf_drainvec_vld[i] ? ibuf_dual : (ibuf_byp & ldst_dual_r) & (i == WrPtr1_r));
			assign buf_dualtag_in[i * DEPTH_LOG2+:DEPTH_LOG2] = (ibuf_drainvec_vld[i] ? ibuf_dualtag : ((ibuf_byp & ldst_dual_r) & (i == WrPtr1_r) ? WrPtr0_r : WrPtr1_r));
			assign buf_sideeffect_in[i] = (ibuf_drainvec_vld[i] ? ibuf_sideeffect : is_sideeffects_r);
			assign buf_unsign_in[i] = (ibuf_drainvec_vld[i] ? ibuf_unsign : lsu_pkt_r[5]);
			assign buf_sz_in[i * 2+:2] = (ibuf_drainvec_vld[i] ? ibuf_sz : {lsu_pkt_r[9], lsu_pkt_r[10]});
			assign buf_write_in[i] = (ibuf_drainvec_vld[i] ? ibuf_write : lsu_pkt_r[6]);
			function automatic [DEPTH_LOG2 - 1:0] sv2v_cast_63A9F;
				input reg [DEPTH_LOG2 - 1:0] inp;
				sv2v_cast_63A9F = inp;
			endfunction
			function automatic signed [pt[181-:8] - 1:0] sv2v_cast_72B45_signed;
				input reg signed [pt[181-:8] - 1:0] inp;
				sv2v_cast_72B45_signed = inp;
			endfunction
			function automatic [pt[181-:8] - 1:0] sv2v_cast_72B45;
				input reg [pt[181-:8] - 1:0] inp;
				sv2v_cast_72B45 = inp;
			endfunction
			function automatic signed [DEPTH_LOG2 - 1:0] sv2v_cast_63A9F_signed;
				input reg signed [DEPTH_LOG2 - 1:0] inp;
				sv2v_cast_63A9F_signed = inp;
			endfunction
			always @(*) begin
				buf_nxtstate[i * 3+:3] = IDLE;
				buf_state_en[i] = 1'b0;
				buf_resp_state_bus_en[i] = 1'b0;
				buf_state_bus_en[i] = 1'b0;
				buf_wr_en[i] = 1'b0;
				buf_data_in[i * 32+:32] = {32 {1'sb0}};
				buf_data_en[i] = 1'b0;
				buf_error_en[i] = 1'b0;
				buf_rst[i] = dec_tlu_force_halt;
				buf_ldfwd_en[i] = dec_tlu_force_halt;
				buf_ldfwd_in[i] = 1'b0;
				buf_ldfwdtag_in[i * DEPTH_LOG2+:DEPTH_LOG2] = {DEPTH_LOG2 {1'sb0}};
				case (buf_state[i * 3+:3])
					IDLE: begin
						buf_nxtstate[i * 3+:3] = (lsu_bus_clk_en ? CMD : WAIT);
						buf_state_en[i] = ((lsu_busreq_r & lsu_commit_r) & ((((ibuf_byp | ldst_dual_r) & ~ibuf_merge_en) & (i == WrPtr0_r)) | ((ibuf_byp & ldst_dual_r) & (i == WrPtr1_r)))) | (ibuf_drain_vld & (i == ibuf_tag));
						buf_wr_en[i] = buf_state_en[i];
						buf_data_en[i] = buf_state_en[i];
						buf_data_in[i * 32+:32] = (ibuf_drain_vld & (i == ibuf_tag) ? ibuf_data_out[31:0] : store_data_lo_r[31:0]);
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					WAIT: begin
						buf_nxtstate[i * 3+:3] = (dec_tlu_force_halt ? IDLE : CMD);
						buf_state_en[i] = lsu_bus_clk_en | dec_tlu_force_halt;
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					CMD: begin
						buf_nxtstate[i * 3+:3] = (dec_tlu_force_halt ? IDLE : ((obuf_nosend & bus_rsp_read) & (bus_rsp_read_tag == obuf_rdrsp_tag) ? DONE_WAIT : RESP));
						buf_cmd_state_bus_en[i] = (((obuf_tag0 == i) | (obuf_merge & (obuf_tag1 == i))) & obuf_valid) & obuf_wr_enQ;
						buf_state_bus_en[i] = buf_cmd_state_bus_en[i];
						buf_state_en[i] = (buf_state_bus_en[i] & lsu_bus_clk_en) | dec_tlu_force_halt;
						buf_ldfwd_in[i] = 1'b1;
						buf_ldfwd_en[i] = ((buf_state_en[i] & ~buf_write[i]) & obuf_nosend) & ~dec_tlu_force_halt;
						buf_ldfwdtag_in[i * DEPTH_LOG2+:DEPTH_LOG2] = sv2v_cast_63A9F(obuf_rdrsp_tag[pt[181-:8] - 2:0]);
						buf_data_en[i] = ((buf_state_bus_en[i] & lsu_bus_clk_en) & obuf_nosend) & bus_rsp_read;
						buf_error_en[i] = ((buf_state_bus_en[i] & lsu_bus_clk_en) & obuf_nosend) & bus_rsp_read_error;
						buf_data_in[i * 32+:32] = (buf_error_en[i] ? bus_rsp_rdata[31:0] : (buf_addr[(i * 32) + 2] ? bus_rsp_rdata[63:32] : bus_rsp_rdata[31:0]));
					end
					RESP: begin
						buf_nxtstate[i * 3+:3] = (dec_tlu_force_halt | (buf_write[i] & ~bus_rsp_write_error) ? IDLE : (((buf_dual[i] & ~buf_samedw[i]) & ~buf_write[i]) & (buf_state[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2] * 3+:3] != DONE_PARTIAL) ? DONE_PARTIAL : ((buf_ldfwd[i] | any_done_wait_state) | (((((buf_dual[i] & ~buf_samedw[i]) & ~buf_write[i]) & buf_ldfwd[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2]]) & (buf_state[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2] * 3+:3] == DONE_PARTIAL)) & any_done_wait_state) ? DONE_WAIT : DONE)));
						buf_resp_state_bus_en[i] = (bus_rsp_write & (bus_rsp_write_tag == sv2v_cast_72B45_signed(i))) | (bus_rsp_read & (((bus_rsp_read_tag == sv2v_cast_72B45_signed(i)) | (buf_ldfwd[i] & (bus_rsp_read_tag == sv2v_cast_72B45(buf_ldfwdtag[i * DEPTH_LOG2+:DEPTH_LOG2])))) | ((((buf_dual[i] & buf_dualhi[i]) & ~buf_write[i]) & buf_samedw[i]) & (bus_rsp_read_tag == sv2v_cast_72B45(buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2])))));
						buf_state_bus_en[i] = buf_resp_state_bus_en[i];
						buf_state_en[i] = (buf_state_bus_en[i] & lsu_bus_clk_en) | dec_tlu_force_halt;
						buf_data_en[i] = (buf_state_bus_en[i] & bus_rsp_read) & lsu_bus_clk_en;
						buf_error_en[i] = (buf_state_bus_en[i] & lsu_bus_clk_en) & (((bus_rsp_read_error & (bus_rsp_read_tag == sv2v_cast_72B45_signed(i))) | ((bus_rsp_read_error & buf_ldfwd[i]) & (bus_rsp_read_tag == sv2v_cast_72B45(buf_ldfwdtag[i * DEPTH_LOG2+:DEPTH_LOG2])))) | (bus_rsp_write_error & (bus_rsp_write_tag == sv2v_cast_72B45_signed(i))));
						buf_data_in[(i * 32) + 31-:32] = (buf_state_en[i] & ~buf_error_en[i] ? (buf_addr[(i * 32) + 2] ? bus_rsp_rdata[63:32] : bus_rsp_rdata[31:0]) : bus_rsp_rdata[31:0]);
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					DONE_PARTIAL: begin
						buf_nxtstate[i * 3+:3] = (dec_tlu_force_halt ? IDLE : ((buf_ldfwd[i] | buf_ldfwd[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2]]) | any_done_wait_state ? DONE_WAIT : DONE));
						buf_state_bus_en[i] = bus_rsp_read & ((bus_rsp_read_tag == sv2v_cast_72B45(buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2])) | (buf_ldfwd[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2]] & (bus_rsp_read_tag == sv2v_cast_72B45(buf_ldfwdtag[buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2] * DEPTH_LOG2+:DEPTH_LOG2]))));
						buf_state_en[i] = (buf_state_bus_en[i] & lsu_bus_clk_en) | dec_tlu_force_halt;
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					DONE_WAIT: begin
						buf_nxtstate[i * 3+:3] = (dec_tlu_force_halt ? IDLE : DONE);
						buf_state_en[i] = ((RspPtr == sv2v_cast_63A9F_signed(i)) | (buf_dual[i] & (buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2] == RspPtr))) | dec_tlu_force_halt;
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					DONE: begin
						buf_nxtstate[i * 3+:3] = IDLE;
						buf_rst[i] = 1'b1;
						buf_state_en[i] = 1'b1;
						buf_ldfwd_in[i] = 1'b0;
						buf_ldfwd_en[i] = buf_state_en[i];
						buf_cmd_state_bus_en[i] = 1'b0;
					end
					default: begin
						buf_nxtstate[i * 3+:3] = IDLE;
						buf_state_en[i] = 1'b0;
						buf_resp_state_bus_en[i] = 1'b0;
						buf_state_bus_en[i] = 1'b0;
						buf_wr_en[i] = 1'b0;
						buf_data_in[i * 32+:32] = {32 {1'sb0}};
						buf_data_en[i] = 1'b0;
						buf_error_en[i] = 1'b0;
						buf_rst[i] = 1'b0;
						buf_cmd_state_bus_en[i] = 1'b0;
					end
				endcase
			end
			rvdffs #(.WIDTH(3)) buf_state_ff(
				.din(buf_nxtstate[i * 3+:3]),
				.dout({buf_state[i * 3+:3]}),
				.en(buf_state_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(DEPTH)) buf_ageff(
				.din(buf_age_in[i * DEPTH+:DEPTH]),
				.dout(buf_ageQ[i * DEPTH+:DEPTH]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(DEPTH)) buf_rspageff(
				.din(buf_rspage_in[i * DEPTH+:DEPTH]),
				.dout(buf_rspageQ[i * DEPTH+:DEPTH]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(DEPTH_LOG2)) buf_dualtagff(
				.din(buf_dualtag_in[i * DEPTH_LOG2+:DEPTH_LOG2]),
				.dout(buf_dualtag[i * DEPTH_LOG2+:DEPTH_LOG2]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_dualff(
				.din(buf_dual_in[i]),
				.dout(buf_dual[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_samedwff(
				.din(buf_samedw_in[i]),
				.dout(buf_samedw[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_nomergeff(
				.din(buf_nomerge_in[i]),
				.dout(buf_nomerge[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_dualhiff(
				.din(buf_dualhi_in[i]),
				.dout(buf_dualhi[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_ldfwdff(
				.din(buf_ldfwd_in[i]),
				.dout(buf_ldfwd[i]),
				.en(buf_ldfwd_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(DEPTH_LOG2)) buf_ldfwdtagff(
				.din(buf_ldfwdtag_in[i * DEPTH_LOG2+:DEPTH_LOG2]),
				.dout(buf_ldfwdtag[i * DEPTH_LOG2+:DEPTH_LOG2]),
				.en(buf_ldfwd_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_sideeffectff(
				.din(buf_sideeffect_in[i]),
				.dout(buf_sideeffect[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_unsignff(
				.din(buf_unsign_in[i]),
				.dout(buf_unsign[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(1)) buf_writeff(
				.din(buf_write_in[i]),
				.dout(buf_write[i]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffs #(.WIDTH(2)) buf_szff(
				.din(buf_sz_in[i * 2+:2]),
				.dout(buf_sz[i * 2+:2]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffe #(.WIDTH(32)) buf_addrff(
				.din(buf_addr_in[(i * 32) + 31-:32]),
				.dout(buf_addr[i * 32+:32]),
				.en(buf_wr_en[i]),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
			rvdffs #(.WIDTH(4)) buf_byteenff(
				.din(buf_byteen_in[(i * 4) + 3-:4]),
				.dout(buf_byteen[i * 4+:4]),
				.en(buf_wr_en[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
			rvdffe #(.WIDTH(32)) buf_dataff(
				.din(buf_data_in[(i * 32) + 31-:32]),
				.dout(buf_data[i * 32+:32]),
				.en(buf_data_en[i]),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
			rvdffsc #(.WIDTH(1)) buf_errorff(
				.din(1'b1),
				.dout(buf_error[i]),
				.en(buf_error_en[i]),
				.clear(buf_rst[i]),
				.clk(lsu_bus_buf_c1_clk),
				.rst_l(rst_l)
			);
		end
	endgenerate
	always @(*) begin
		buf_numvld_any[3:0] = (({1'b0, lsu_busreq_m} << ldst_dual_m) + ({1'b0, lsu_busreq_r} << ldst_dual_r)) + ibuf_valid;
		buf_numvld_wrcmd_any[3:0] = 4'b0000;
		buf_numvld_cmd_any[3:0] = 4'b0000;
		buf_numvld_pend_any[3:0] = 4'b0000;
		any_done_wait_state = 1'b0;
		begin : sv2v_autoblock_53
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					buf_numvld_any[3:0] = buf_numvld_any[3:0] + {3'b000, buf_state[i * 3+:3] != IDLE};
					buf_numvld_wrcmd_any[3:0] = buf_numvld_wrcmd_any[3:0] + {3'b000, (buf_write[i] & (buf_state[i * 3+:3] == CMD)) & ~buf_cmd_state_bus_en[i]};
					buf_numvld_cmd_any[3:0] = buf_numvld_cmd_any[3:0] + {3'b000, (buf_state[i * 3+:3] == CMD) & ~buf_cmd_state_bus_en[i]};
					buf_numvld_pend_any[3:0] = buf_numvld_pend_any[3:0] + {3'b000, (buf_state[i * 3+:3] == WAIT) | ((buf_state[i * 3+:3] == CMD) & ~buf_cmd_state_bus_en[i])};
					any_done_wait_state = any_done_wait_state | (buf_state[i * 3+:3] == DONE_WAIT);
				end
		end
	end
	assign lsu_bus_buffer_pend_any = buf_numvld_pend_any != 0;
	assign lsu_bus_buffer_full_any = (ldst_dual_d & dec_lsu_valid_raw_d ? buf_numvld_any[3:0] >= (DEPTH - 1) : buf_numvld_any[3:0] == DEPTH);
	assign lsu_bus_buffer_empty_any = (~(|buf_state[3 * ((DEPTH - 1) - (DEPTH - 1))+:3 * DEPTH]) & ~ibuf_valid) & ~obuf_valid;
	assign lsu_nonblock_load_valid_m = (((lsu_busreq_m & lsu_pkt_m[0]) & lsu_pkt_m[7]) & ~flush_m_up) & ~ld_full_hit_m;
	assign lsu_nonblock_load_tag_m[DEPTH_LOG2 - 1:0] = WrPtr0_m[DEPTH_LOG2 - 1:0];
	assign lsu_nonblock_load_inv_r = lsu_nonblock_load_valid_r & ~lsu_commit_r;
	assign lsu_nonblock_load_inv_tag_r[DEPTH_LOG2 - 1:0] = WrPtr0_r[DEPTH_LOG2 - 1:0];
	always @(*) begin
		lsu_nonblock_load_data_ready = 1'b0;
		lsu_nonblock_load_data_error = 1'b0;
		lsu_nonblock_load_data_tag[DEPTH_LOG2 - 1:0] = {DEPTH_LOG2 {1'sb0}};
		lsu_nonblock_load_data_lo[31:0] = {32 {1'sb0}};
		lsu_nonblock_load_data_hi[31:0] = {32 {1'sb0}};
		begin : sv2v_autoblock_54
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					lsu_nonblock_load_data_ready = lsu_nonblock_load_data_ready | ((buf_state[i * 3+:3] == DONE) & ~buf_write[i]);
					lsu_nonblock_load_data_error = lsu_nonblock_load_data_error | (((buf_state[i * 3+:3] == DONE) & buf_error[i]) & ~buf_write[i]);
					lsu_nonblock_load_data_tag[DEPTH_LOG2 - 1:0] = lsu_nonblock_load_data_tag[DEPTH_LOG2 - 1:0] | (sv2v_cast_63A9F_signed(i) & {DEPTH_LOG2 {((buf_state[i * 3+:3] == DONE) & ~buf_write[i]) & (~buf_dual[i] | ~buf_dualhi[i])}});
					lsu_nonblock_load_data_lo[31:0] = lsu_nonblock_load_data_lo[31:0] | (buf_data[(i * 32) + 31-:32] & {32 {((buf_state[i * 3+:3] == DONE) & ~buf_write[i]) & (~buf_dual[i] | ~buf_dualhi[i])}});
					lsu_nonblock_load_data_hi[31:0] = lsu_nonblock_load_data_hi[31:0] | (buf_data[(i * 32) + 31-:32] & {32 {((buf_state[i * 3+:3] == DONE) & ~buf_write[i]) & (buf_dual[i] & buf_dualhi[i])}});
				end
		end
	end
	assign lsu_nonblock_addr_offset[1:0] = buf_addr[(lsu_nonblock_load_data_tag * 32) + 1-:2];
	assign lsu_nonblock_sz[1:0] = buf_sz[(lsu_nonblock_load_data_tag * 2) + 1-:2];
	assign lsu_nonblock_unsign = buf_unsign[lsu_nonblock_load_data_tag];
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign lsu_nonblock_data_unalgn[31:0] = sv2v_cast_32({lsu_nonblock_load_data_hi[31:0], lsu_nonblock_load_data_lo[31:0]} >> (8 * lsu_nonblock_addr_offset[1:0]));
	assign lsu_nonblock_load_data_valid = lsu_nonblock_load_data_ready & ~lsu_nonblock_load_data_error;
	assign lsu_nonblock_load_data[31:0] = (((({32 {lsu_nonblock_unsign & (lsu_nonblock_sz[1:0] == 2'b00)}} & {24'b000000000000000000000000, lsu_nonblock_data_unalgn[7:0]}) | ({32 {lsu_nonblock_unsign & (lsu_nonblock_sz[1:0] == 2'b01)}} & {16'b0000000000000000, lsu_nonblock_data_unalgn[15:0]})) | ({32 {~lsu_nonblock_unsign & (lsu_nonblock_sz[1:0] == 2'b00)}} & {{24 {lsu_nonblock_data_unalgn[7]}}, lsu_nonblock_data_unalgn[7:0]})) | ({32 {~lsu_nonblock_unsign & (lsu_nonblock_sz[1:0] == 2'b01)}} & {{16 {lsu_nonblock_data_unalgn[15]}}, lsu_nonblock_data_unalgn[15:0]})) | ({32 {lsu_nonblock_sz[1:0] == 2'b10}} & lsu_nonblock_data_unalgn[31:0]);
	always @(*) begin
		bus_sideeffect_pend = (obuf_valid & obuf_sideeffect) & dec_tlu_sideeffect_posted_disable;
		begin : sv2v_autoblock_55
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				bus_sideeffect_pend = bus_sideeffect_pend | (((buf_state[i * 3+:3] == RESP) & buf_sideeffect[i]) & dec_tlu_sideeffect_posted_disable);
		end
	end
	function automatic signed [pt[181-:8] - 1:0] sv2v_cast_72B45_signed;
		input reg signed [pt[181-:8] - 1:0] inp;
		sv2v_cast_72B45_signed = inp;
	endfunction
	always @(*) begin
		bus_addr_match_pending = 1'b0;
		begin : sv2v_autoblock_56
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				bus_addr_match_pending = bus_addr_match_pending | (((obuf_valid & (obuf_addr[31:3] == buf_addr[(i * 32) + 31-:29])) & (buf_state[i * 3+:3] == RESP)) & ~((obuf_tag0 == sv2v_cast_72B45_signed(i)) | (obuf_merge & (obuf_tag1 == sv2v_cast_72B45_signed(i)))));
		end
	end
	assign bus_cmd_ready = (obuf_write ? (obuf_cmd_done | obuf_data_done ? (obuf_cmd_done ? lsu_axi_wready : lsu_axi_awready) : lsu_axi_awready & lsu_axi_wready) : lsu_axi_arready);
	assign bus_wcmd_sent = lsu_axi_awvalid & lsu_axi_awready;
	assign bus_wdata_sent = lsu_axi_wvalid & lsu_axi_wready;
	assign bus_cmd_sent = ((obuf_cmd_done | bus_wcmd_sent) & (obuf_data_done | bus_wdata_sent)) | (lsu_axi_arvalid & lsu_axi_arready);
	assign bus_rsp_read = lsu_axi_rvalid & lsu_axi_rready;
	assign bus_rsp_write = lsu_axi_bvalid & lsu_axi_bready;
	assign bus_rsp_read_tag[pt[181-:8] - 1:0] = lsu_axi_rid[pt[181-:8] - 1:0];
	assign bus_rsp_write_tag[pt[181-:8] - 1:0] = lsu_axi_bid[pt[181-:8] - 1:0];
	assign bus_rsp_write_error = bus_rsp_write & (lsu_axi_bresp[1:0] != 2'b00);
	assign bus_rsp_read_error = bus_rsp_read & (lsu_axi_rresp[1:0] != 2'b00);
	assign bus_rsp_rdata[63:0] = lsu_axi_rdata[63:0];
	assign lsu_axi_awvalid = ((obuf_valid & obuf_write) & ~obuf_cmd_done) & ~bus_addr_match_pending;
	assign lsu_axi_awid[pt[181-:8] - 1:0] = sv2v_cast_72B45(obuf_tag0);
	assign lsu_axi_awaddr[31:0] = (obuf_sideeffect ? obuf_addr[31:0] : {obuf_addr[31:3], 3'b000});
	assign lsu_axi_awsize[2:0] = (obuf_sideeffect ? {1'b0, obuf_sz[1:0]} : 3'b011);
	assign lsu_axi_awprot[2:0] = 3'b001;
	assign lsu_axi_awcache[3:0] = (obuf_sideeffect ? 4'b0000 : 4'b1111);
	assign lsu_axi_awregion[3:0] = obuf_addr[31:28];
	assign lsu_axi_awlen[7:0] = {8 {1'sb0}};
	assign lsu_axi_awburst[1:0] = 2'b01;
	assign lsu_axi_awqos[3:0] = {4 {1'sb0}};
	assign lsu_axi_awlock = 1'b0;
	assign lsu_axi_wvalid = ((obuf_valid & obuf_write) & ~obuf_data_done) & ~bus_addr_match_pending;
	assign lsu_axi_wstrb[7:0] = obuf_byteen[7:0] & {8 {obuf_write}};
	assign lsu_axi_wdata[63:0] = obuf_data[63:0];
	assign lsu_axi_wlast = 1'b1;
	assign lsu_axi_arvalid = ((obuf_valid & ~obuf_write) & ~obuf_nosend) & ~bus_addr_match_pending;
	assign lsu_axi_arid[pt[181-:8] - 1:0] = sv2v_cast_72B45(obuf_tag0);
	assign lsu_axi_araddr[31:0] = (obuf_sideeffect ? obuf_addr[31:0] : {obuf_addr[31:3], 3'b000});
	assign lsu_axi_arsize[2:0] = (obuf_sideeffect ? {1'b0, obuf_sz[1:0]} : 3'b011);
	assign lsu_axi_arprot[2:0] = 3'b001;
	assign lsu_axi_arcache[3:0] = (obuf_sideeffect ? 4'b0000 : 4'b1111);
	assign lsu_axi_arregion[3:0] = obuf_addr[31:28];
	assign lsu_axi_arlen[7:0] = {8 {1'sb0}};
	assign lsu_axi_arburst[1:0] = 2'b01;
	assign lsu_axi_arqos[3:0] = {4 {1'sb0}};
	assign lsu_axi_arlock = 1'b0;
	assign lsu_axi_bready = 1;
	assign lsu_axi_rready = 1;
	always @(*) begin
		lsu_imprecise_error_store_any = 1'b0;
		lsu_imprecise_error_store_tag = {pt[181-:8] {1'sb0}};
		begin : sv2v_autoblock_57
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					lsu_imprecise_error_store_any = lsu_imprecise_error_store_any | (((lsu_bus_clk_en_q & (buf_state[i * 3+:3] == DONE)) & buf_error[i]) & buf_write[i]);
					lsu_imprecise_error_store_tag = lsu_imprecise_error_store_tag | (sv2v_cast_63A9F_signed(i) & {DEPTH_LOG2 {((buf_state[i * 3+:3] == DONE) & buf_error[i]) & buf_write[i]}});
				end
		end
	end
	assign lsu_imprecise_error_load_any = lsu_nonblock_load_data_error & ~lsu_imprecise_error_store_any;
	assign lsu_imprecise_error_addr_any[31:0] = (lsu_imprecise_error_store_any ? buf_addr[lsu_imprecise_error_store_tag * 32+:32] : buf_addr[lsu_nonblock_load_data_tag * 32+:32]);
	assign lsu_pmu_bus_trxn = ((lsu_axi_awvalid & lsu_axi_awready) | (lsu_axi_wvalid & lsu_axi_wready)) | (lsu_axi_arvalid & lsu_axi_arready);
	assign lsu_pmu_bus_misaligned = (lsu_busreq_r & ldst_dual_r) & lsu_commit_r;
	assign lsu_pmu_bus_error = lsu_imprecise_error_load_any | lsu_imprecise_error_store_any;
	assign lsu_pmu_bus_busy = ((lsu_axi_awvalid & ~lsu_axi_awready) | (lsu_axi_wvalid & ~lsu_axi_wready)) | (lsu_axi_arvalid & ~lsu_axi_arready);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_awvalid_ff(
		.din(lsu_axi_awvalid),
		.dout(lsu_axi_awvalid_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_awready_ff(
		.din(lsu_axi_awready),
		.dout(lsu_axi_awready_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_wvalid_ff(
		.din(lsu_axi_wvalid),
		.dout(lsu_axi_wvalid_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_wready_ff(
		.din(lsu_axi_wready),
		.dout(lsu_axi_wready_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_arvalid_ff(
		.din(lsu_axi_arvalid),
		.dout(lsu_axi_arvalid_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_arready_ff(
		.din(lsu_axi_arready),
		.dout(lsu_axi_arready_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_bvalid_ff(
		.din(lsu_axi_bvalid),
		.dout(lsu_axi_bvalid_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_bready_ff(
		.din(lsu_axi_bready),
		.dout(lsu_axi_bready_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(2)) lsu_axi_bresp_ff(
		.din(lsu_axi_bresp[1:0]),
		.dout(lsu_axi_bresp_q[1:0]),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(pt[181-:8])) lsu_axi_bid_ff(
		.din(lsu_axi_bid[pt[181-:8] - 1:0]),
		.dout(lsu_axi_bid_q[pt[181-:8] - 1:0]),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(64)) lsu_axi_rdata_ff(
		.din(lsu_axi_rdata[63:0]),
		.dout(lsu_axi_rdata_q[63:0]),
		.en((lsu_axi_rvalid | clk_override) & lsu_bus_clk_en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_rvalid_ff(
		.din(lsu_axi_rvalid),
		.dout(lsu_axi_rvalid_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(1)) lsu_axi_rready_ff(
		.din(lsu_axi_rready),
		.dout(lsu_axi_rready_q),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(2)) lsu_axi_rresp_ff(
		.din(lsu_axi_rresp[1:0]),
		.dout(lsu_axi_rresp_q[1:0]),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff_fpga #(.WIDTH(pt[181-:8])) lsu_axi_rid_ff(
		.din(lsu_axi_rid[pt[181-:8] - 1:0]),
		.dout(lsu_axi_rid_q[pt[181-:8] - 1:0]),
		.clk(lsu_busm_clk),
		.clken(lsu_busm_clken),
		.rawclk(clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(DEPTH_LOG2)) lsu_WrPtr0_rff(
		.din(WrPtr0_m),
		.dout(WrPtr0_r),
		.clk(lsu_c2_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(DEPTH_LOG2)) lsu_WrPtr1_rff(
		.din(WrPtr1_m),
		.dout(WrPtr1_r),
		.clk(lsu_c2_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) lsu_busreq_rff(
		.din((lsu_busreq_m & ~flush_r) & ~ld_full_hit_m),
		.dout(lsu_busreq_r),
		.clk(lsu_c2_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) lsu_nonblock_load_valid_rff(
		.din(lsu_nonblock_load_valid_m),
		.dout(lsu_nonblock_load_valid_r),
		.clk(lsu_c2_r_clk),
		.rst_l(rst_l)
	);
endmodule
module eb1_lsu_bus_intf (
	clk,
	clk_override,
	rst_l,
	scan_mode,
	dec_tlu_external_ldfwd_disable,
	dec_tlu_wb_coalescing_disable,
	dec_tlu_sideeffect_posted_disable,
	lsu_bus_obuf_c1_clken,
	lsu_busm_clken,
	lsu_c1_r_clk,
	lsu_c2_r_clk,
	lsu_bus_ibuf_c1_clk,
	lsu_bus_obuf_c1_clk,
	lsu_bus_buf_c1_clk,
	lsu_free_c2_clk,
	active_clk,
	lsu_busm_clk,
	dec_lsu_valid_raw_d,
	lsu_busreq_m,
	lsu_pkt_m,
	lsu_pkt_r,
	lsu_addr_m,
	lsu_addr_r,
	end_addr_m,
	end_addr_r,
	store_data_r,
	dec_tlu_force_halt,
	lsu_commit_r,
	is_sideeffects_m,
	flush_m_up,
	flush_r,
	ldst_dual_d,
	ldst_dual_m,
	ldst_dual_r,
	lsu_busreq_r,
	lsu_bus_buffer_pend_any,
	lsu_bus_buffer_full_any,
	lsu_bus_buffer_empty_any,
	bus_read_data_m,
	lsu_imprecise_error_load_any,
	lsu_imprecise_error_store_any,
	lsu_imprecise_error_addr_any,
	lsu_nonblock_load_valid_m,
	lsu_nonblock_load_tag_m,
	lsu_nonblock_load_inv_r,
	lsu_nonblock_load_inv_tag_r,
	lsu_nonblock_load_data_valid,
	lsu_nonblock_load_data_error,
	lsu_nonblock_load_data_tag,
	lsu_nonblock_load_data,
	lsu_pmu_bus_trxn,
	lsu_pmu_bus_misaligned,
	lsu_pmu_bus_error,
	lsu_pmu_bus_busy,
	lsu_axi_awvalid,
	lsu_axi_awready,
	lsu_axi_awid,
	lsu_axi_awaddr,
	lsu_axi_awregion,
	lsu_axi_awlen,
	lsu_axi_awsize,
	lsu_axi_awburst,
	lsu_axi_awlock,
	lsu_axi_awcache,
	lsu_axi_awprot,
	lsu_axi_awqos,
	lsu_axi_wvalid,
	lsu_axi_wready,
	lsu_axi_wdata,
	lsu_axi_wstrb,
	lsu_axi_wlast,
	lsu_axi_bvalid,
	lsu_axi_bready,
	lsu_axi_bresp,
	lsu_axi_bid,
	lsu_axi_arvalid,
	lsu_axi_arready,
	lsu_axi_arid,
	lsu_axi_araddr,
	lsu_axi_arregion,
	lsu_axi_arlen,
	lsu_axi_arsize,
	lsu_axi_arburst,
	lsu_axi_arlock,
	lsu_axi_arcache,
	lsu_axi_arprot,
	lsu_axi_arqos,
	lsu_axi_rvalid,
	lsu_axi_rready,
	lsu_axi_rid,
	lsu_axi_rdata,
	lsu_axi_rresp,
	lsu_bus_clk_en
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire clk_override;
	input wire rst_l;
	input wire scan_mode;
	input wire dec_tlu_external_ldfwd_disable;
	input wire dec_tlu_wb_coalescing_disable;
	input wire dec_tlu_sideeffect_posted_disable;
	input wire lsu_bus_obuf_c1_clken;
	input wire lsu_busm_clken;
	input wire lsu_c1_r_clk;
	input wire lsu_c2_r_clk;
	input wire lsu_bus_ibuf_c1_clk;
	input wire lsu_bus_obuf_c1_clk;
	input wire lsu_bus_buf_c1_clk;
	input wire lsu_free_c2_clk;
	input wire active_clk;
	input wire lsu_busm_clk;
	input wire dec_lsu_valid_raw_d;
	input wire lsu_busreq_m;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_r;
	input wire [31:0] lsu_addr_m;
	input wire [31:0] lsu_addr_r;
	input wire [31:0] end_addr_m;
	input wire [31:0] end_addr_r;
	input wire [31:0] store_data_r;
	input wire dec_tlu_force_halt;
	input wire lsu_commit_r;
	input wire is_sideeffects_m;
	input wire flush_m_up;
	input wire flush_r;
	input wire ldst_dual_d;
	input wire ldst_dual_m;
	input wire ldst_dual_r;
	output wire lsu_busreq_r;
	output wire lsu_bus_buffer_pend_any;
	output wire lsu_bus_buffer_full_any;
	output wire lsu_bus_buffer_empty_any;
	output wire [31:0] bus_read_data_m;
	output wire lsu_imprecise_error_load_any;
	output wire lsu_imprecise_error_store_any;
	output wire [31:0] lsu_imprecise_error_addr_any;
	output wire lsu_nonblock_load_valid_m;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_tag_m;
	output wire lsu_nonblock_load_inv_r;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_inv_tag_r;
	output wire lsu_nonblock_load_data_valid;
	output wire lsu_nonblock_load_data_error;
	output wire [pt[164-:7] - 1:0] lsu_nonblock_load_data_tag;
	output wire [31:0] lsu_nonblock_load_data;
	output wire lsu_pmu_bus_trxn;
	output wire lsu_pmu_bus_misaligned;
	output wire lsu_pmu_bus_error;
	output wire lsu_pmu_bus_busy;
	output wire lsu_axi_awvalid;
	input wire lsu_axi_awready;
	output wire [pt[181-:8] - 1:0] lsu_axi_awid;
	output wire [31:0] lsu_axi_awaddr;
	output wire [3:0] lsu_axi_awregion;
	output wire [7:0] lsu_axi_awlen;
	output wire [2:0] lsu_axi_awsize;
	output wire [1:0] lsu_axi_awburst;
	output wire lsu_axi_awlock;
	output wire [3:0] lsu_axi_awcache;
	output wire [2:0] lsu_axi_awprot;
	output wire [3:0] lsu_axi_awqos;
	output wire lsu_axi_wvalid;
	input wire lsu_axi_wready;
	output wire [63:0] lsu_axi_wdata;
	output wire [7:0] lsu_axi_wstrb;
	output wire lsu_axi_wlast;
	input wire lsu_axi_bvalid;
	output wire lsu_axi_bready;
	input wire [1:0] lsu_axi_bresp;
	input wire [pt[181-:8] - 1:0] lsu_axi_bid;
	output wire lsu_axi_arvalid;
	input wire lsu_axi_arready;
	output wire [pt[181-:8] - 1:0] lsu_axi_arid;
	output wire [31:0] lsu_axi_araddr;
	output wire [3:0] lsu_axi_arregion;
	output wire [7:0] lsu_axi_arlen;
	output wire [2:0] lsu_axi_arsize;
	output wire [1:0] lsu_axi_arburst;
	output wire lsu_axi_arlock;
	output wire [3:0] lsu_axi_arcache;
	output wire [2:0] lsu_axi_arprot;
	output wire [3:0] lsu_axi_arqos;
	input wire lsu_axi_rvalid;
	output wire lsu_axi_rready;
	input wire [pt[181-:8] - 1:0] lsu_axi_rid;
	input wire [63:0] lsu_axi_rdata;
	input wire [1:0] lsu_axi_rresp;
	input wire lsu_bus_clk_en;
	wire lsu_bus_clk_en_q;
	wire [3:0] ldst_byteen_m;
	wire [3:0] ldst_byteen_r;
	wire [7:0] ldst_byteen_ext_m;
	wire [7:0] ldst_byteen_ext_r;
	wire [3:0] ldst_byteen_hi_m;
	wire [3:0] ldst_byteen_hi_r;
	wire [3:0] ldst_byteen_lo_m;
	wire [3:0] ldst_byteen_lo_r;
	wire is_sideeffects_r;
	wire [63:0] store_data_ext_r;
	wire [31:0] store_data_hi_r;
	wire [31:0] store_data_lo_r;
	wire addr_match_dw_lo_r_m;
	wire addr_match_word_lo_r_m;
	wire no_word_merge_r;
	wire no_dword_merge_r;
	wire ld_addr_rhit_lo_lo;
	wire ld_addr_rhit_hi_lo;
	wire ld_addr_rhit_lo_hi;
	wire ld_addr_rhit_hi_hi;
	wire [3:0] ld_byte_rhit_lo_lo;
	wire [3:0] ld_byte_rhit_hi_lo;
	wire [3:0] ld_byte_rhit_lo_hi;
	wire [3:0] ld_byte_rhit_hi_hi;
	wire [3:0] ld_byte_hit_lo;
	wire [3:0] ld_byte_rhit_lo;
	wire [3:0] ld_byte_hit_hi;
	wire [3:0] ld_byte_rhit_hi;
	wire [31:0] ld_fwddata_rpipe_lo;
	wire [31:0] ld_fwddata_rpipe_hi;
	wire [3:0] ld_byte_hit_buf_lo;
	wire [3:0] ld_byte_hit_buf_hi;
	wire [31:0] ld_fwddata_buf_lo;
	wire [31:0] ld_fwddata_buf_hi;
	wire [63:0] ld_fwddata_lo;
	wire [63:0] ld_fwddata_hi;
	wire [63:0] ld_fwddata_m;
	reg ld_full_hit_hi_m;
	reg ld_full_hit_lo_m;
	wire ld_full_hit_m;
	assign ldst_byteen_m[3:0] = (({4 {lsu_pkt_m[11]}} & 4'b0001) | ({4 {lsu_pkt_m[10]}} & 4'b0011)) | ({4 {lsu_pkt_m[9]}} & 4'b1111);
	eb1_lsu_bus_buffer #(.pt(pt)) bus_buffer(
		.clk(clk),
		.clk_override(clk_override),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.dec_tlu_external_ldfwd_disable(dec_tlu_external_ldfwd_disable),
		.dec_tlu_wb_coalescing_disable(dec_tlu_wb_coalescing_disable),
		.dec_tlu_sideeffect_posted_disable(dec_tlu_sideeffect_posted_disable),
		.dec_tlu_force_halt(dec_tlu_force_halt),
		.lsu_bus_obuf_c1_clken(lsu_bus_obuf_c1_clken),
		.lsu_busm_clken(lsu_busm_clken),
		.lsu_c2_r_clk(lsu_c2_r_clk),
		.lsu_bus_ibuf_c1_clk(lsu_bus_ibuf_c1_clk),
		.lsu_bus_obuf_c1_clk(lsu_bus_obuf_c1_clk),
		.lsu_bus_buf_c1_clk(lsu_bus_buf_c1_clk),
		.lsu_free_c2_clk(lsu_free_c2_clk),
		.lsu_busm_clk(lsu_busm_clk),
		.dec_lsu_valid_raw_d(dec_lsu_valid_raw_d),
		.lsu_pkt_m(lsu_pkt_m),
		.lsu_pkt_r(lsu_pkt_r),
		.lsu_addr_m(lsu_addr_m),
		.end_addr_m(end_addr_m),
		.lsu_addr_r(lsu_addr_r),
		.end_addr_r(end_addr_r),
		.store_data_r(store_data_r),
		.no_word_merge_r(no_word_merge_r),
		.no_dword_merge_r(no_dword_merge_r),
		.lsu_busreq_m(lsu_busreq_m),
		.lsu_busreq_r(lsu_busreq_r),
		.ld_full_hit_m(ld_full_hit_m),
		.flush_m_up(flush_m_up),
		.flush_r(flush_r),
		.lsu_commit_r(lsu_commit_r),
		.is_sideeffects_r(is_sideeffects_r),
		.ldst_dual_d(ldst_dual_d),
		.ldst_dual_m(ldst_dual_m),
		.ldst_dual_r(ldst_dual_r),
		.ldst_byteen_ext_m(ldst_byteen_ext_m),
		.lsu_bus_buffer_pend_any(lsu_bus_buffer_pend_any),
		.lsu_bus_buffer_full_any(lsu_bus_buffer_full_any),
		.lsu_bus_buffer_empty_any(lsu_bus_buffer_empty_any),
		.ld_byte_hit_buf_lo(ld_byte_hit_buf_lo),
		.ld_byte_hit_buf_hi(ld_byte_hit_buf_hi),
		.ld_fwddata_buf_lo(ld_fwddata_buf_lo),
		.ld_fwddata_buf_hi(ld_fwddata_buf_hi),
		.lsu_imprecise_error_load_any(lsu_imprecise_error_load_any),
		.lsu_imprecise_error_store_any(lsu_imprecise_error_store_any),
		.lsu_imprecise_error_addr_any(lsu_imprecise_error_addr_any),
		.lsu_nonblock_load_valid_m(lsu_nonblock_load_valid_m),
		.lsu_nonblock_load_tag_m(lsu_nonblock_load_tag_m),
		.lsu_nonblock_load_inv_r(lsu_nonblock_load_inv_r),
		.lsu_nonblock_load_inv_tag_r(lsu_nonblock_load_inv_tag_r),
		.lsu_nonblock_load_data_valid(lsu_nonblock_load_data_valid),
		.lsu_nonblock_load_data_error(lsu_nonblock_load_data_error),
		.lsu_nonblock_load_data_tag(lsu_nonblock_load_data_tag),
		.lsu_nonblock_load_data(lsu_nonblock_load_data),
		.lsu_pmu_bus_trxn(lsu_pmu_bus_trxn),
		.lsu_pmu_bus_misaligned(lsu_pmu_bus_misaligned),
		.lsu_pmu_bus_error(lsu_pmu_bus_error),
		.lsu_pmu_bus_busy(lsu_pmu_bus_busy),
		.lsu_axi_awvalid(lsu_axi_awvalid),
		.lsu_axi_awready(lsu_axi_awready),
		.lsu_axi_awid(lsu_axi_awid),
		.lsu_axi_awaddr(lsu_axi_awaddr),
		.lsu_axi_awregion(lsu_axi_awregion),
		.lsu_axi_awlen(lsu_axi_awlen),
		.lsu_axi_awsize(lsu_axi_awsize),
		.lsu_axi_awburst(lsu_axi_awburst),
		.lsu_axi_awlock(lsu_axi_awlock),
		.lsu_axi_awcache(lsu_axi_awcache),
		.lsu_axi_awprot(lsu_axi_awprot),
		.lsu_axi_awqos(lsu_axi_awqos),
		.lsu_axi_wvalid(lsu_axi_wvalid),
		.lsu_axi_wready(lsu_axi_wready),
		.lsu_axi_wdata(lsu_axi_wdata),
		.lsu_axi_wstrb(lsu_axi_wstrb),
		.lsu_axi_wlast(lsu_axi_wlast),
		.lsu_axi_bvalid(lsu_axi_bvalid),
		.lsu_axi_bready(lsu_axi_bready),
		.lsu_axi_bresp(lsu_axi_bresp),
		.lsu_axi_bid(lsu_axi_bid),
		.lsu_axi_arvalid(lsu_axi_arvalid),
		.lsu_axi_arready(lsu_axi_arready),
		.lsu_axi_arid(lsu_axi_arid),
		.lsu_axi_araddr(lsu_axi_araddr),
		.lsu_axi_arregion(lsu_axi_arregion),
		.lsu_axi_arlen(lsu_axi_arlen),
		.lsu_axi_arsize(lsu_axi_arsize),
		.lsu_axi_arburst(lsu_axi_arburst),
		.lsu_axi_arlock(lsu_axi_arlock),
		.lsu_axi_arcache(lsu_axi_arcache),
		.lsu_axi_arprot(lsu_axi_arprot),
		.lsu_axi_arqos(lsu_axi_arqos),
		.lsu_axi_rvalid(lsu_axi_rvalid),
		.lsu_axi_rready(lsu_axi_rready),
		.lsu_axi_rid(lsu_axi_rid),
		.lsu_axi_rdata(lsu_axi_rdata),
		.lsu_axi_rresp(lsu_axi_rresp),
		.lsu_bus_clk_en(lsu_bus_clk_en),
		.lsu_bus_clk_en_q(lsu_bus_clk_en_q)
	);
	assign addr_match_dw_lo_r_m = lsu_addr_r[31:3] == lsu_addr_m[31:3];
	assign addr_match_word_lo_r_m = addr_match_dw_lo_r_m & ~(lsu_addr_r[2] ^ lsu_addr_m[2]);
	assign no_word_merge_r = ((lsu_busreq_r & ~ldst_dual_r) & lsu_busreq_m) & (lsu_pkt_m[7] | ~addr_match_word_lo_r_m);
	assign no_dword_merge_r = ((lsu_busreq_r & ~ldst_dual_r) & lsu_busreq_m) & (lsu_pkt_m[7] | ~addr_match_dw_lo_r_m);
	assign ldst_byteen_ext_m[7:0] = {4'b0000, ldst_byteen_m[3:0]} << lsu_addr_m[1:0];
	assign ldst_byteen_ext_r[7:0] = {4'b0000, ldst_byteen_r[3:0]} << lsu_addr_r[1:0];
	assign store_data_ext_r[63:0] = {32'b00000000000000000000000000000000, store_data_r[31:0]} << {lsu_addr_r[1:0], 3'b000};
	assign ldst_byteen_hi_m[3:0] = ldst_byteen_ext_m[7:4];
	assign ldst_byteen_lo_m[3:0] = ldst_byteen_ext_m[3:0];
	assign ldst_byteen_hi_r[3:0] = ldst_byteen_ext_r[7:4];
	assign ldst_byteen_lo_r[3:0] = ldst_byteen_ext_r[3:0];
	assign store_data_hi_r[31:0] = store_data_ext_r[63:32];
	assign store_data_lo_r[31:0] = store_data_ext_r[31:0];
	assign ld_addr_rhit_lo_lo = (((lsu_addr_m[31:2] == lsu_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & lsu_busreq_m;
	assign ld_addr_rhit_lo_hi = (((end_addr_m[31:2] == lsu_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & lsu_busreq_m;
	assign ld_addr_rhit_hi_lo = (((lsu_addr_m[31:2] == end_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & lsu_busreq_m;
	assign ld_addr_rhit_hi_hi = (((end_addr_m[31:2] == end_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & lsu_busreq_m;
	generate
		genvar i;
		for (i = 0; i < 4; i = i + 1) begin : GenBusBufFwd
			assign ld_byte_rhit_lo_lo[i] = (ld_addr_rhit_lo_lo & ldst_byteen_lo_r[i]) & ldst_byteen_lo_m[i];
			assign ld_byte_rhit_lo_hi[i] = (ld_addr_rhit_lo_hi & ldst_byteen_lo_r[i]) & ldst_byteen_hi_m[i];
			assign ld_byte_rhit_hi_lo[i] = (ld_addr_rhit_hi_lo & ldst_byteen_hi_r[i]) & ldst_byteen_lo_m[i];
			assign ld_byte_rhit_hi_hi[i] = (ld_addr_rhit_hi_hi & ldst_byteen_hi_r[i]) & ldst_byteen_hi_m[i];
			assign ld_byte_hit_lo[i] = (ld_byte_rhit_lo_lo[i] | ld_byte_rhit_hi_lo[i]) | ld_byte_hit_buf_lo[i];
			assign ld_byte_hit_hi[i] = (ld_byte_rhit_lo_hi[i] | ld_byte_rhit_hi_hi[i]) | ld_byte_hit_buf_hi[i];
			assign ld_byte_rhit_lo[i] = ld_byte_rhit_lo_lo[i] | ld_byte_rhit_hi_lo[i];
			assign ld_byte_rhit_hi[i] = ld_byte_rhit_lo_hi[i] | ld_byte_rhit_hi_hi[i];
			assign ld_fwddata_rpipe_lo[(8 * i) + 7:8 * i] = ({8 {ld_byte_rhit_lo_lo[i]}} & store_data_lo_r[(8 * i) + 7:8 * i]) | ({8 {ld_byte_rhit_hi_lo[i]}} & store_data_hi_r[(8 * i) + 7:8 * i]);
			assign ld_fwddata_rpipe_hi[(8 * i) + 7:8 * i] = ({8 {ld_byte_rhit_lo_hi[i]}} & store_data_lo_r[(8 * i) + 7:8 * i]) | ({8 {ld_byte_rhit_hi_hi[i]}} & store_data_hi_r[(8 * i) + 7:8 * i]);
			assign ld_fwddata_lo[(8 * i) + 7:8 * i] = (ld_byte_rhit_lo[i] ? ld_fwddata_rpipe_lo[(8 * i) + 7:8 * i] : ld_fwddata_buf_lo[(8 * i) + 7:8 * i]);
			assign ld_fwddata_hi[(8 * i) + 7:8 * i] = (ld_byte_rhit_hi[i] ? ld_fwddata_rpipe_hi[(8 * i) + 7:8 * i] : ld_fwddata_buf_hi[(8 * i) + 7:8 * i]);
		end
	endgenerate
	always @(*) begin
		ld_full_hit_lo_m = 1'b1;
		ld_full_hit_hi_m = 1'b1;
		begin : sv2v_autoblock_58
			reg signed [31:0] i;
			for (i = 0; i < 4; i = i + 1)
				begin
					ld_full_hit_lo_m = ld_full_hit_lo_m & (ld_byte_hit_lo[i] | ~ldst_byteen_lo_m[i]);
					ld_full_hit_hi_m = ld_full_hit_hi_m & (ld_byte_hit_hi[i] | ~ldst_byteen_hi_m[i]);
				end
		end
	end
	assign ld_full_hit_m = (((ld_full_hit_lo_m & ld_full_hit_hi_m) & lsu_busreq_m) & lsu_pkt_m[7]) & ~is_sideeffects_m;
	assign ld_fwddata_m[63:0] = {ld_fwddata_hi[31:0], ld_fwddata_lo[31:0]} >> (8 * lsu_addr_m[1:0]);
	assign bus_read_data_m[31:0] = ld_fwddata_m[31:0];
	rvdff #(.WIDTH(1)) clken_ff(
		.din(lsu_bus_clk_en),
		.dout(lsu_bus_clk_en_q),
		.clk(active_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) is_sideeffects_rff(
		.din(is_sideeffects_m),
		.dout(is_sideeffects_r),
		.clk(lsu_c1_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(4)) lsu_byten_rff(
		.rst_l(rst_l),
		.din(ldst_byteen_m[3:0]),
		.dout(ldst_byteen_r[3:0]),
		.clk(lsu_c1_r_clk)
	);
endmodule
module eb1_lsu_clkdomain (
	clk,
	active_clk,
	rst_l,
	dec_tlu_force_halt,
	clk_override,
	dma_dccm_req,
	ldst_stbuf_reqvld_r,
	stbuf_reqvld_any,
	stbuf_reqvld_flushed_any,
	lsu_busreq_r,
	lsu_bus_buffer_pend_any,
	lsu_bus_buffer_empty_any,
	lsu_stbuf_empty_any,
	lsu_bus_clk_en,
	lsu_p,
	lsu_pkt_d,
	lsu_pkt_m,
	lsu_pkt_r,
	lsu_bus_obuf_c1_clken,
	lsu_busm_clken,
	lsu_c1_m_clk,
	lsu_c1_r_clk,
	lsu_c2_m_clk,
	lsu_c2_r_clk,
	lsu_store_c1_m_clk,
	lsu_store_c1_r_clk,
	lsu_stbuf_c1_clk,
	lsu_bus_obuf_c1_clk,
	lsu_bus_ibuf_c1_clk,
	lsu_bus_buf_c1_clk,
	lsu_busm_clk,
	lsu_free_c2_clk,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire active_clk;
	input wire rst_l;
	input wire dec_tlu_force_halt;
	input wire clk_override;
	input wire dma_dccm_req;
	input wire ldst_stbuf_reqvld_r;
	input wire stbuf_reqvld_any;
	input wire stbuf_reqvld_flushed_any;
	input wire lsu_busreq_r;
	input wire lsu_bus_buffer_pend_any;
	input wire lsu_bus_buffer_empty_any;
	input wire lsu_stbuf_empty_any;
	input wire lsu_bus_clk_en;
	input wire [13:0] lsu_p;
	input wire [13:0] lsu_pkt_d;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_r;
	output wire lsu_bus_obuf_c1_clken;
	output wire lsu_busm_clken;
	output wire lsu_c1_m_clk;
	output wire lsu_c1_r_clk;
	output wire lsu_c2_m_clk;
	output wire lsu_c2_r_clk;
	output wire lsu_store_c1_m_clk;
	output wire lsu_store_c1_r_clk;
	output wire lsu_stbuf_c1_clk;
	output wire lsu_bus_obuf_c1_clk;
	output wire lsu_bus_ibuf_c1_clk;
	output wire lsu_bus_buf_c1_clk;
	output wire lsu_busm_clk;
	output wire lsu_free_c2_clk;
	input wire scan_mode;
	wire lsu_c1_m_clken;
	wire lsu_c1_r_clken;
	wire lsu_c2_m_clken;
	wire lsu_c2_r_clken;
	wire lsu_c1_m_clken_q;
	wire lsu_c1_r_clken_q;
	wire lsu_store_c1_m_clken;
	wire lsu_store_c1_r_clken;
	wire lsu_stbuf_c1_clken;
	wire lsu_bus_ibuf_c1_clken;
	wire lsu_bus_buf_c1_clken;
	wire lsu_free_c1_clken;
	wire lsu_free_c1_clken_q;
	wire lsu_free_c2_clken;
	assign lsu_c1_m_clken = (lsu_p[0] | dma_dccm_req) | clk_override;
	assign lsu_c1_r_clken = (lsu_pkt_m[0] | lsu_c1_m_clken_q) | clk_override;
	assign lsu_c2_m_clken = (lsu_c1_m_clken | lsu_c1_m_clken_q) | clk_override;
	assign lsu_c2_r_clken = (lsu_c1_r_clken | lsu_c1_r_clken_q) | clk_override;
	assign lsu_store_c1_m_clken = (lsu_c1_m_clken & lsu_pkt_d[6]) | clk_override;
	assign lsu_store_c1_r_clken = (lsu_c1_r_clken & lsu_pkt_m[6]) | clk_override;
	assign lsu_stbuf_c1_clken = ((ldst_stbuf_reqvld_r | stbuf_reqvld_any) | stbuf_reqvld_flushed_any) | clk_override;
	assign lsu_bus_ibuf_c1_clken = lsu_busreq_r | clk_override;
	assign lsu_bus_obuf_c1_clken = ((lsu_bus_buffer_pend_any | lsu_busreq_r) | clk_override) & lsu_bus_clk_en;
	assign lsu_bus_buf_c1_clken = ((~lsu_bus_buffer_empty_any | lsu_busreq_r) | dec_tlu_force_halt) | clk_override;
	assign lsu_free_c1_clken = (((((lsu_p[0] | lsu_pkt_d[0]) | lsu_pkt_m[0]) | lsu_pkt_r[0]) | ~lsu_bus_buffer_empty_any) | ~lsu_stbuf_empty_any) | clk_override;
	assign lsu_free_c2_clken = (lsu_free_c1_clken | lsu_free_c1_clken_q) | clk_override;
	rvdff #(.WIDTH(1)) lsu_free_c1_clkenff(
		.din(lsu_free_c1_clken),
		.dout(lsu_free_c1_clken_q),
		.clk(active_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) lsu_c1_m_clkenff(
		.din(lsu_c1_m_clken),
		.dout(lsu_c1_m_clken_q),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) lsu_c1_r_clkenff(
		.din(lsu_c1_r_clken),
		.dout(lsu_c1_r_clken_q),
		.clk(lsu_free_c2_clk),
		.rst_l(rst_l)
	);
	rvoclkhdr lsu_c1m_cgc(
		.en(lsu_c1_m_clken),
		.l1clk(lsu_c1_m_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_c1r_cgc(
		.en(lsu_c1_r_clken),
		.l1clk(lsu_c1_r_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_c2m_cgc(
		.en(lsu_c2_m_clken),
		.l1clk(lsu_c2_m_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_c2r_cgc(
		.en(lsu_c2_r_clken),
		.l1clk(lsu_c2_r_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_store_c1m_cgc(
		.en(lsu_store_c1_m_clken),
		.l1clk(lsu_store_c1_m_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_store_c1r_cgc(
		.en(lsu_store_c1_r_clken),
		.l1clk(lsu_store_c1_r_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_stbuf_c1_cgc(
		.en(lsu_stbuf_c1_clken),
		.l1clk(lsu_stbuf_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_bus_ibuf_c1_cgc(
		.en(lsu_bus_ibuf_c1_clken),
		.l1clk(lsu_bus_ibuf_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_bus_buf_c1_cgc(
		.en(lsu_bus_buf_c1_clken),
		.l1clk(lsu_bus_buf_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	assign lsu_busm_clken = ((~lsu_bus_buffer_empty_any | lsu_busreq_r) | clk_override) & lsu_bus_clk_en;
	rvclkhdr lsu_bus_obuf_c1_cgc(
		.en(lsu_bus_obuf_c1_clken),
		.l1clk(lsu_bus_obuf_c1_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvclkhdr lsu_busm_cgc(
		.en(lsu_busm_clken),
		.l1clk(lsu_busm_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
	rvoclkhdr lsu_free_cgc(
		.en(lsu_free_c2_clken),
		.l1clk(lsu_free_c2_clk),
		.clk(clk),
		.scan_mode(scan_mode)
	);
endmodule
module eb1_lsu_dccm_ctl (
	lsu_c2_m_clk,
	lsu_c2_r_clk,
	lsu_c1_r_clk,
	lsu_store_c1_r_clk,
	lsu_free_c2_clk,
	clk_override,
	clk,
	rst_l,
	lsu_pkt_r,
	lsu_pkt_m,
	lsu_pkt_d,
	addr_in_dccm_d,
	addr_in_pic_d,
	addr_in_pic_m,
	addr_in_dccm_m,
	addr_in_dccm_r,
	addr_in_pic_r,
	lsu_raw_fwd_lo_r,
	lsu_raw_fwd_hi_r,
	lsu_commit_r,
	ldst_dual_m,
	ldst_dual_r,
	lsu_addr_d,
	lsu_addr_m,
	lsu_addr_r,
	end_addr_d,
	end_addr_m,
	end_addr_r,
	stbuf_reqvld_any,
	stbuf_addr_any,
	stbuf_data_any,
	stbuf_ecc_any,
	stbuf_fwddata_hi_m,
	stbuf_fwddata_lo_m,
	stbuf_fwdbyteen_hi_m,
	stbuf_fwdbyteen_lo_m,
	dccm_rdata_hi_r,
	dccm_rdata_lo_r,
	dccm_data_ecc_hi_r,
	dccm_data_ecc_lo_r,
	lsu_ld_data_r,
	lsu_ld_data_corr_r,
	lsu_double_ecc_error_r,
	single_ecc_error_hi_r,
	single_ecc_error_lo_r,
	sec_data_hi_r,
	sec_data_lo_r,
	sec_data_hi_r_ff,
	sec_data_lo_r_ff,
	sec_data_ecc_hi_r_ff,
	sec_data_ecc_lo_r_ff,
	dccm_rdata_hi_m,
	dccm_rdata_lo_m,
	dccm_data_ecc_hi_m,
	dccm_data_ecc_lo_m,
	lsu_ld_data_m,
	lsu_double_ecc_error_m,
	sec_data_hi_m,
	sec_data_lo_m,
	store_data_m,
	dma_dccm_wen,
	dma_pic_wen,
	dma_mem_tag_m,
	dma_mem_addr,
	dma_mem_wdata,
	dma_dccm_wdata_lo,
	dma_dccm_wdata_hi,
	dma_dccm_wdata_ecc_hi,
	dma_dccm_wdata_ecc_lo,
	store_data_hi_r,
	store_data_lo_r,
	store_datafn_hi_r,
	store_datafn_lo_r,
	store_data_r,
	ld_single_ecc_error_r,
	ld_single_ecc_error_r_ff,
	picm_mask_data_m,
	lsu_stbuf_commit_any,
	lsu_dccm_rden_m,
	lsu_dccm_rden_r,
	dccm_dma_rvalid,
	dccm_dma_ecc_error,
	dccm_dma_rtag,
	dccm_dma_rdata,
	dccm_wren,
	dccm_rden,
	dccm_wr_addr_lo,
	dccm_wr_addr_hi,
	dccm_rd_addr_lo,
	dccm_rd_addr_hi,
	dccm_wr_data_lo,
	dccm_wr_data_hi,
	dccm_rd_data_lo,
	dccm_rd_data_hi,
	picm_wren,
	picm_rden,
	picm_mken,
	picm_rdaddr,
	picm_wraddr,
	picm_wr_data,
	picm_rd_data,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire lsu_c2_m_clk;
	input wire lsu_c2_r_clk;
	input wire lsu_c1_r_clk;
	input wire lsu_store_c1_r_clk;
	input wire lsu_free_c2_clk;
	input wire clk_override;
	input wire clk;
	input wire rst_l;
	input wire [13:0] lsu_pkt_r;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_d;
	input wire addr_in_dccm_d;
	input wire addr_in_pic_d;
	input wire addr_in_pic_m;
	input wire addr_in_dccm_m;
	input wire addr_in_dccm_r;
	input wire addr_in_pic_r;
	input wire lsu_raw_fwd_lo_r;
	input wire lsu_raw_fwd_hi_r;
	input wire lsu_commit_r;
	input wire ldst_dual_m;
	input wire ldst_dual_r;
	input wire [31:0] lsu_addr_d;
	input wire [pt[1398-:9] - 1:0] lsu_addr_m;
	input wire [31:0] lsu_addr_r;
	input wire [pt[1398-:9] - 1:0] end_addr_d;
	input wire [pt[1398-:9] - 1:0] end_addr_m;
	input wire [pt[1398-:9] - 1:0] end_addr_r;
	input wire stbuf_reqvld_any;
	input wire [pt[157-:9] - 1:0] stbuf_addr_any;
	input wire [pt[1382-:10] - 1:0] stbuf_data_any;
	input wire [pt[1372-:7] - 1:0] stbuf_ecc_any;
	input wire [pt[1382-:10] - 1:0] stbuf_fwddata_hi_m;
	input wire [pt[1382-:10] - 1:0] stbuf_fwddata_lo_m;
	input wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_hi_m;
	input wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_lo_m;
	output wire [pt[1382-:10] - 1:0] dccm_rdata_hi_r;
	output wire [pt[1382-:10] - 1:0] dccm_rdata_lo_r;
	output wire [pt[1372-:7] - 1:0] dccm_data_ecc_hi_r;
	output wire [pt[1372-:7] - 1:0] dccm_data_ecc_lo_r;
	output wire [pt[1382-:10] - 1:0] lsu_ld_data_r;
	output wire [pt[1382-:10] - 1:0] lsu_ld_data_corr_r;
	input wire lsu_double_ecc_error_r;
	input wire single_ecc_error_hi_r;
	input wire single_ecc_error_lo_r;
	input wire [pt[1382-:10] - 1:0] sec_data_hi_r;
	input wire [pt[1382-:10] - 1:0] sec_data_lo_r;
	input wire [pt[1382-:10] - 1:0] sec_data_hi_r_ff;
	input wire [pt[1382-:10] - 1:0] sec_data_lo_r_ff;
	input wire [pt[1372-:7] - 1:0] sec_data_ecc_hi_r_ff;
	input wire [pt[1372-:7] - 1:0] sec_data_ecc_lo_r_ff;
	output wire [pt[1382-:10] - 1:0] dccm_rdata_hi_m;
	output wire [pt[1382-:10] - 1:0] dccm_rdata_lo_m;
	output wire [pt[1372-:7] - 1:0] dccm_data_ecc_hi_m;
	output wire [pt[1372-:7] - 1:0] dccm_data_ecc_lo_m;
	output wire [pt[1382-:10] - 1:0] lsu_ld_data_m;
	input wire lsu_double_ecc_error_m;
	input wire [pt[1382-:10] - 1:0] sec_data_hi_m;
	input wire [pt[1382-:10] - 1:0] sec_data_lo_m;
	input wire [31:0] store_data_m;
	input wire dma_dccm_wen;
	input wire dma_pic_wen;
	input wire [2:0] dma_mem_tag_m;
	input wire [31:0] dma_mem_addr;
	input wire [63:0] dma_mem_wdata;
	input wire [31:0] dma_dccm_wdata_lo;
	input wire [31:0] dma_dccm_wdata_hi;
	input wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_hi;
	input wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_lo;
	output wire [pt[1382-:10] - 1:0] store_data_hi_r;
	output wire [pt[1382-:10] - 1:0] store_data_lo_r;
	output wire [pt[1382-:10] - 1:0] store_datafn_hi_r;
	output wire [pt[1382-:10] - 1:0] store_datafn_lo_r;
	output wire [31:0] store_data_r;
	output wire ld_single_ecc_error_r;
	output wire ld_single_ecc_error_r_ff;
	output wire [31:0] picm_mask_data_m;
	output wire lsu_stbuf_commit_any;
	output wire lsu_dccm_rden_m;
	output wire lsu_dccm_rden_r;
	output wire dccm_dma_rvalid;
	output wire dccm_dma_ecc_error;
	output wire [2:0] dccm_dma_rtag;
	output wire [63:0] dccm_dma_rdata;
	output wire dccm_wren;
	output wire dccm_rden;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	output wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	output wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	input wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	output wire picm_wren;
	output wire picm_rden;
	output wire picm_mken;
	output wire [31:0] picm_rdaddr;
	output wire [31:0] picm_wraddr;
	output wire [31:0] picm_wr_data;
	input wire [31:0] picm_rd_data;
	input wire scan_mode;
	localparam DCCM_WIDTH_BITS = $clog2(pt[1389-:7]);
	wire lsu_dccm_rden_d;
	wire lsu_dccm_wren_d;
	wire ld_single_ecc_error_lo_r;
	wire ld_single_ecc_error_hi_r;
	wire ld_single_ecc_error_lo_r_ns;
	wire ld_single_ecc_error_hi_r_ns;
	wire ld_single_ecc_error_lo_r_ff;
	wire ld_single_ecc_error_hi_r_ff;
	wire lsu_double_ecc_error_r_ff;
	wire [pt[1398-:9] - 1:0] ld_sec_addr_lo_r_ff;
	wire [pt[1398-:9] - 1:0] ld_sec_addr_hi_r_ff;
	wire [pt[1382-:10] - 1:0] store_data_lo_r_in;
	wire [pt[1382-:10] - 1:0] store_data_hi_r_in;
	wire [63:0] picm_rd_data_m;
	wire dccm_wr_bypass_d_m_hi;
	wire dccm_wr_bypass_d_r_hi;
	wire dccm_wr_bypass_d_m_lo;
	wire dccm_wr_bypass_d_r_lo;
	wire kill_ecc_corr_lo_r;
	wire kill_ecc_corr_hi_r;
	wire [3:0] store_byteen_m;
	wire [3:0] store_byteen_r;
	wire [7:0] store_byteen_ext_m;
	wire [7:0] store_byteen_ext_r;
	generate
		if (pt[202-:5] == 1) begin : L2U_Plus1_1
			wire [63:0] lsu_rdata_r;
			wire [63:0] lsu_rdata_corr_r;
			wire [63:0] dccm_rdata_r;
			wire [63:0] dccm_rdata_corr_r;
			wire [63:0] stbuf_fwddata_r;
			wire [7:0] stbuf_fwdbyteen_r;
			wire [31:0] stbuf_fwddata_lo_r;
			wire [31:0] stbuf_fwddata_hi_r;
			wire [3:0] stbuf_fwdbyteen_lo_r;
			wire [3:0] stbuf_fwdbyteen_hi_r;
			wire [31:0] lsu_rdata_lo_r;
			wire [31:0] lsu_rdata_hi_r;
			wire [63:0] picm_rd_data_r;
			wire [63:32] lsu_ld_data_r_nc;
			wire [63:32] lsu_ld_data_corr_r_nc;
			wire [2:0] dma_mem_tag_r;
			wire stbuf_fwddata_en;
			assign dccm_dma_rvalid = (lsu_pkt_r[0] & lsu_pkt_r[7]) & lsu_pkt_r[4];
			assign dccm_dma_ecc_error = lsu_double_ecc_error_r;
			assign dccm_dma_rtag[2:0] = dma_mem_tag_r[2:0];
			assign dccm_dma_rdata[63:0] = (ldst_dual_r ? lsu_rdata_corr_r[63:0] : {2 {lsu_rdata_corr_r[31:0]}});
			assign {lsu_ld_data_r_nc[63:32], lsu_ld_data_r[31:0]} = lsu_rdata_r[63:0] >> (8 * lsu_addr_r[1:0]);
			assign {lsu_ld_data_corr_r_nc[63:32], lsu_ld_data_corr_r[31:0]} = lsu_rdata_corr_r[63:0] >> (8 * lsu_addr_r[1:0]);
			assign picm_rd_data_r[63:32] = picm_rd_data_r[31:0];
			assign dccm_rdata_r[63:0] = {dccm_rdata_hi_r[31:0], dccm_rdata_lo_r[31:0]};
			assign dccm_rdata_corr_r[63:0] = {sec_data_hi_r[31:0], sec_data_lo_r[31:0]};
			assign stbuf_fwddata_r[63:0] = {stbuf_fwddata_hi_r[31:0], stbuf_fwddata_lo_r[31:0]};
			assign stbuf_fwdbyteen_r[7:0] = {stbuf_fwdbyteen_hi_r[3:0], stbuf_fwdbyteen_lo_r[3:0]};
			assign stbuf_fwddata_en = (|stbuf_fwdbyteen_hi_m[3:0] | |stbuf_fwdbyteen_lo_m[3:0]) | clk_override;
			genvar i;
			for (i = 0; i < 8; i = i + 1) begin : GenDMAData
				assign lsu_rdata_corr_r[(8 * i) + 7:8 * i] = (stbuf_fwdbyteen_r[i] ? stbuf_fwddata_r[(8 * i) + 7:8 * i] : (addr_in_pic_r ? picm_rd_data_r[(8 * i) + 7:8 * i] : {8 {addr_in_dccm_r}} & dccm_rdata_corr_r[(8 * i) + 7:8 * i]));
				assign lsu_rdata_r[(8 * i) + 7:8 * i] = (stbuf_fwdbyteen_r[i] ? stbuf_fwddata_r[(8 * i) + 7:8 * i] : (addr_in_pic_r ? picm_rd_data_r[(8 * i) + 7:8 * i] : {8 {addr_in_dccm_r}} & dccm_rdata_r[(8 * i) + 7:8 * i]));
			end
			rvdffe #(.WIDTH(pt[1382-:10])) dccm_rdata_hi_r_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(dccm_rdata_hi_m[pt[1382-:10] - 1:0]),
				.dout(dccm_rdata_hi_r[pt[1382-:10] - 1:0]),
				.en((lsu_dccm_rden_m & ldst_dual_m) | clk_override)
			);
			rvdffe #(.WIDTH(pt[1382-:10])) dccm_rdata_lo_r_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(dccm_rdata_lo_m[pt[1382-:10] - 1:0]),
				.dout(dccm_rdata_lo_r[pt[1382-:10] - 1:0]),
				.en(lsu_dccm_rden_m | clk_override)
			);
			rvdffe #(.WIDTH(2 * pt[1372-:7])) dccm_data_ecc_r_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din({dccm_data_ecc_hi_m[pt[1372-:7] - 1:0], dccm_data_ecc_lo_m[pt[1372-:7] - 1:0]}),
				.dout({dccm_data_ecc_hi_r[pt[1372-:7] - 1:0], dccm_data_ecc_lo_r[pt[1372-:7] - 1:0]}),
				.en(lsu_dccm_rden_m | clk_override)
			);
			rvdff #(.WIDTH(8)) stbuf_fwdbyteen_ff(
				.rst_l(rst_l),
				.din({stbuf_fwdbyteen_hi_m[3:0], stbuf_fwdbyteen_lo_m[3:0]}),
				.dout({stbuf_fwdbyteen_hi_r[3:0], stbuf_fwdbyteen_lo_r[3:0]}),
				.clk(lsu_c2_r_clk)
			);
			rvdffe #(.WIDTH(64)) stbuf_fwddata_ff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din({stbuf_fwddata_hi_m[31:0], stbuf_fwddata_lo_m[31:0]}),
				.dout({stbuf_fwddata_hi_r[31:0], stbuf_fwddata_lo_r[31:0]}),
				.en(stbuf_fwddata_en)
			);
			rvdffe #(.WIDTH(32)) picm_rddata_rff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(picm_rd_data_m[31:0]),
				.dout(picm_rd_data_r[31:0]),
				.en(addr_in_pic_m | clk_override)
			);
			rvdff #(.WIDTH(3)) dma_mem_tag_rff(
				.rst_l(rst_l),
				.din(dma_mem_tag_m[2:0]),
				.dout(dma_mem_tag_r[2:0]),
				.clk(lsu_c1_r_clk)
			);
		end
		else begin : L2U_Plus1_0
			wire [63:0] lsu_rdata_m;
			wire [63:0] lsu_rdata_corr_m;
			wire [63:0] dccm_rdata_m;
			wire [63:0] dccm_rdata_corr_m;
			wire [63:0] stbuf_fwddata_m;
			wire [7:0] stbuf_fwdbyteen_m;
			wire [63:32] lsu_ld_data_m_nc;
			wire [63:32] lsu_ld_data_corr_m_nc;
			wire [31:0] lsu_ld_data_corr_m;
			assign dccm_dma_rvalid = (lsu_pkt_m[0] & lsu_pkt_m[7]) & lsu_pkt_m[4];
			assign dccm_dma_ecc_error = lsu_double_ecc_error_m;
			assign dccm_dma_rtag[2:0] = dma_mem_tag_m[2:0];
			assign dccm_dma_rdata[63:0] = (ldst_dual_m ? lsu_rdata_corr_m[63:0] : {2 {lsu_rdata_corr_m[31:0]}});
			assign {lsu_ld_data_m_nc[63:32], lsu_ld_data_m[31:0]} = lsu_rdata_m[63:0] >> (8 * lsu_addr_m[1:0]);
			assign {lsu_ld_data_corr_m_nc[63:32], lsu_ld_data_corr_m[31:0]} = lsu_rdata_corr_m[63:0] >> (8 * lsu_addr_m[1:0]);
			assign dccm_rdata_m[63:0] = {dccm_rdata_hi_m[31:0], dccm_rdata_lo_m[31:0]};
			assign dccm_rdata_corr_m[63:0] = {sec_data_hi_m[31:0], sec_data_lo_m[31:0]};
			assign stbuf_fwddata_m[63:0] = {stbuf_fwddata_hi_m[31:0], stbuf_fwddata_lo_m[31:0]};
			assign stbuf_fwdbyteen_m[7:0] = {stbuf_fwdbyteen_hi_m[3:0], stbuf_fwdbyteen_lo_m[3:0]};
			genvar i;
			for (i = 0; i < 8; i = i + 1) begin : GenLoop
				assign lsu_rdata_corr_m[(8 * i) + 7:8 * i] = (stbuf_fwdbyteen_m[i] ? stbuf_fwddata_m[(8 * i) + 7:8 * i] : (addr_in_pic_m ? picm_rd_data_m[(8 * i) + 7:8 * i] : {8 {addr_in_dccm_m}} & dccm_rdata_corr_m[(8 * i) + 7:8 * i]));
				assign lsu_rdata_m[(8 * i) + 7:8 * i] = (stbuf_fwdbyteen_m[i] ? stbuf_fwddata_m[(8 * i) + 7:8 * i] : (addr_in_pic_m ? picm_rd_data_m[(8 * i) + 7:8 * i] : {8 {addr_in_dccm_m}} & dccm_rdata_m[(8 * i) + 7:8 * i]));
			end
			rvdffe #(.WIDTH(32)) lsu_ld_data_corr_rff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(lsu_ld_data_corr_m[31:0]),
				.dout(lsu_ld_data_corr_r[31:0]),
				.en(((lsu_pkt_m[0] & lsu_pkt_m[7]) & (addr_in_pic_m | addr_in_dccm_m)) | clk_override)
			);
		end
	endgenerate
	assign kill_ecc_corr_lo_r = ((((((lsu_addr_d[pt[1398-:9] - 1:2] == lsu_addr_r[pt[1398-:9] - 1:2]) | (end_addr_d[pt[1398-:9] - 1:2] == lsu_addr_r[pt[1398-:9] - 1:2])) & lsu_pkt_d[0]) & lsu_pkt_d[6]) & lsu_pkt_d[4]) & addr_in_dccm_d) | ((((((lsu_addr_m[pt[1398-:9] - 1:2] == lsu_addr_r[pt[1398-:9] - 1:2]) | (end_addr_m[pt[1398-:9] - 1:2] == lsu_addr_r[pt[1398-:9] - 1:2])) & lsu_pkt_m[0]) & lsu_pkt_m[6]) & lsu_pkt_m[4]) & addr_in_dccm_m);
	assign kill_ecc_corr_hi_r = ((((((lsu_addr_d[pt[1398-:9] - 1:2] == end_addr_r[pt[1398-:9] - 1:2]) | (end_addr_d[pt[1398-:9] - 1:2] == end_addr_r[pt[1398-:9] - 1:2])) & lsu_pkt_d[0]) & lsu_pkt_d[6]) & lsu_pkt_d[4]) & addr_in_dccm_d) | ((((((lsu_addr_m[pt[1398-:9] - 1:2] == end_addr_r[pt[1398-:9] - 1:2]) | (end_addr_m[pt[1398-:9] - 1:2] == end_addr_r[pt[1398-:9] - 1:2])) & lsu_pkt_m[0]) & lsu_pkt_m[6]) & lsu_pkt_m[4]) & addr_in_dccm_m);
	assign ld_single_ecc_error_lo_r = (lsu_pkt_r[7] & single_ecc_error_lo_r) & ~lsu_raw_fwd_lo_r;
	assign ld_single_ecc_error_hi_r = (lsu_pkt_r[7] & single_ecc_error_hi_r) & ~lsu_raw_fwd_hi_r;
	assign ld_single_ecc_error_r = (ld_single_ecc_error_lo_r | ld_single_ecc_error_hi_r) & ~lsu_double_ecc_error_r;
	assign ld_single_ecc_error_lo_r_ns = (ld_single_ecc_error_lo_r & (lsu_commit_r | lsu_pkt_r[4])) & ~kill_ecc_corr_lo_r;
	assign ld_single_ecc_error_hi_r_ns = (ld_single_ecc_error_hi_r & (lsu_commit_r | lsu_pkt_r[4])) & ~kill_ecc_corr_hi_r;
	assign ld_single_ecc_error_r_ff = (ld_single_ecc_error_lo_r_ff | ld_single_ecc_error_hi_r_ff) & ~lsu_double_ecc_error_r_ff;
	assign lsu_stbuf_commit_any = stbuf_reqvld_any & (~((lsu_dccm_rden_d | lsu_dccm_wren_d) | ld_single_ecc_error_r_ff) | (lsu_dccm_rden_d & ~((stbuf_addr_any[pt[1275-:6]+:pt[1405-:7]] == lsu_addr_d[pt[1275-:6]+:pt[1405-:7]]) | (stbuf_addr_any[pt[1275-:6]+:pt[1405-:7]] == end_addr_d[pt[1275-:6]+:pt[1405-:7]]))));
	assign lsu_dccm_rden_d = (lsu_pkt_d[0] & (lsu_pkt_d[7] | (lsu_pkt_d[6] & (~(lsu_pkt_d[9] | lsu_pkt_d[8]) | (lsu_addr_d[1:0] != 2'b00))))) & addr_in_dccm_d;
	assign lsu_dccm_wren_d = dma_dccm_wen;
	assign dccm_wren = (lsu_dccm_wren_d | lsu_stbuf_commit_any) | ld_single_ecc_error_r_ff;
	assign dccm_rden = lsu_dccm_rden_d & addr_in_dccm_d;
	assign dccm_wr_addr_lo[pt[1398-:9] - 1:0] = (ld_single_ecc_error_r_ff ? (ld_single_ecc_error_lo_r_ff ? ld_sec_addr_lo_r_ff[pt[1398-:9] - 1:0] : ld_sec_addr_hi_r_ff[pt[1398-:9] - 1:0]) : (lsu_dccm_wren_d ? lsu_addr_d[pt[1398-:9] - 1:0] : stbuf_addr_any[pt[1398-:9] - 1:0]));
	assign dccm_wr_addr_hi[pt[1398-:9] - 1:0] = (ld_single_ecc_error_r_ff ? (ld_single_ecc_error_hi_r_ff ? ld_sec_addr_hi_r_ff[pt[1398-:9] - 1:0] : ld_sec_addr_lo_r_ff[pt[1398-:9] - 1:0]) : (lsu_dccm_wren_d ? end_addr_d[pt[1398-:9] - 1:0] : stbuf_addr_any[pt[1398-:9] - 1:0]));
	assign dccm_rd_addr_lo[pt[1398-:9] - 1:0] = lsu_addr_d[pt[1398-:9] - 1:0];
	assign dccm_rd_addr_hi[pt[1398-:9] - 1:0] = end_addr_d[pt[1398-:9] - 1:0];
	assign dccm_wr_data_lo[pt[1360-:10] - 1:0] = (ld_single_ecc_error_r_ff ? (ld_single_ecc_error_lo_r_ff ? {sec_data_ecc_lo_r_ff[pt[1372-:7] - 1:0], sec_data_lo_r_ff[pt[1382-:10] - 1:0]} : {sec_data_ecc_hi_r_ff[pt[1372-:7] - 1:0], sec_data_hi_r_ff[pt[1382-:10] - 1:0]}) : (dma_dccm_wen ? {dma_dccm_wdata_ecc_lo[pt[1372-:7] - 1:0], dma_dccm_wdata_lo[pt[1382-:10] - 1:0]} : {stbuf_ecc_any[pt[1372-:7] - 1:0], stbuf_data_any[pt[1382-:10] - 1:0]}));
	assign dccm_wr_data_hi[pt[1360-:10] - 1:0] = (ld_single_ecc_error_r_ff ? (ld_single_ecc_error_hi_r_ff ? {sec_data_ecc_hi_r_ff[pt[1372-:7] - 1:0], sec_data_hi_r_ff[pt[1382-:10] - 1:0]} : {sec_data_ecc_lo_r_ff[pt[1372-:7] - 1:0], sec_data_lo_r_ff[pt[1382-:10] - 1:0]}) : (dma_dccm_wen ? {dma_dccm_wdata_ecc_hi[pt[1372-:7] - 1:0], dma_dccm_wdata_hi[pt[1382-:10] - 1:0]} : {stbuf_ecc_any[pt[1372-:7] - 1:0], stbuf_data_any[pt[1382-:10] - 1:0]}));
	assign store_byteen_m[3:0] = {4 {lsu_pkt_m[6]}} & ((({4 {lsu_pkt_m[11]}} & 4'b0001) | ({4 {lsu_pkt_m[10]}} & 4'b0011)) | ({4 {lsu_pkt_m[9]}} & 4'b1111));
	assign store_byteen_r[3:0] = {4 {lsu_pkt_r[6]}} & ((({4 {lsu_pkt_r[11]}} & 4'b0001) | ({4 {lsu_pkt_r[10]}} & 4'b0011)) | ({4 {lsu_pkt_r[9]}} & 4'b1111));
	assign store_byteen_ext_m[7:0] = {4'b0000, store_byteen_m[3:0]} << lsu_addr_m[1:0];
	assign store_byteen_ext_r[7:0] = {4'b0000, store_byteen_r[3:0]} << lsu_addr_r[1:0];
	assign dccm_wr_bypass_d_m_lo = (stbuf_addr_any[pt[1398-:9] - 1:2] == lsu_addr_m[pt[1398-:9] - 1:2]) & addr_in_dccm_m;
	assign dccm_wr_bypass_d_m_hi = (stbuf_addr_any[pt[1398-:9] - 1:2] == end_addr_m[pt[1398-:9] - 1:2]) & addr_in_dccm_m;
	assign dccm_wr_bypass_d_r_lo = (stbuf_addr_any[pt[1398-:9] - 1:2] == lsu_addr_r[pt[1398-:9] - 1:2]) & addr_in_dccm_r;
	assign dccm_wr_bypass_d_r_hi = (stbuf_addr_any[pt[1398-:9] - 1:2] == end_addr_r[pt[1398-:9] - 1:2]) & addr_in_dccm_r;
	generate
		if (pt[202-:5] == 1) begin : L2U1_Plus1_1
			wire dccm_wren_Q;
			wire [31:0] dccm_wr_data_Q;
			wire dccm_wr_bypass_d_m_lo_Q;
			wire dccm_wr_bypass_d_m_hi_Q;
			wire [31:0] store_data_pre_hi_r;
			wire [31:0] store_data_pre_lo_r;
			assign {store_data_pre_hi_r[31:0], store_data_pre_lo_r[31:0]} = {32'b00000000000000000000000000000000, store_data_r[31:0]} << (8 * lsu_addr_r[1:0]);
			genvar i;
			for (i = 0; i < 4; i = i + 1) begin
				assign store_data_lo_r[(8 * i) + 7:8 * i] = (store_byteen_ext_r[i] ? store_data_pre_lo_r[(8 * i) + 7:8 * i] : (dccm_wren_Q & dccm_wr_bypass_d_m_lo_Q ? dccm_wr_data_Q[(8 * i) + 7:8 * i] : sec_data_lo_r[(8 * i) + 7:8 * i]));
				assign store_data_hi_r[(8 * i) + 7:8 * i] = (store_byteen_ext_r[i + 4] ? store_data_pre_hi_r[(8 * i) + 7:8 * i] : (dccm_wren_Q & dccm_wr_bypass_d_m_hi_Q ? dccm_wr_data_Q[(8 * i) + 7:8 * i] : sec_data_hi_r[(8 * i) + 7:8 * i]));
				assign store_datafn_lo_r[(8 * i) + 7:8 * i] = (store_byteen_ext_r[i] ? store_data_pre_lo_r[(8 * i) + 7:8 * i] : (lsu_stbuf_commit_any & dccm_wr_bypass_d_r_lo ? stbuf_data_any[(8 * i) + 7:8 * i] : (dccm_wren_Q & dccm_wr_bypass_d_m_lo_Q ? dccm_wr_data_Q[(8 * i) + 7:8 * i] : sec_data_lo_r[(8 * i) + 7:8 * i])));
				assign store_datafn_hi_r[(8 * i) + 7:8 * i] = (store_byteen_ext_r[i + 4] ? store_data_pre_hi_r[(8 * i) + 7:8 * i] : (lsu_stbuf_commit_any & dccm_wr_bypass_d_r_hi ? stbuf_data_any[(8 * i) + 7:8 * i] : (dccm_wren_Q & dccm_wr_bypass_d_m_hi_Q ? dccm_wr_data_Q[(8 * i) + 7:8 * i] : sec_data_hi_r[(8 * i) + 7:8 * i])));
			end
			rvdff #(.WIDTH(1)) dccm_wren_ff(
				.rst_l(rst_l),
				.din(lsu_stbuf_commit_any),
				.dout(dccm_wren_Q),
				.clk(lsu_free_c2_clk)
			);
			rvdffe #(.WIDTH(32)) dccm_wrdata_ff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(stbuf_data_any[31:0]),
				.dout(dccm_wr_data_Q[31:0]),
				.en(lsu_stbuf_commit_any | clk_override),
				.clk(clk)
			);
			rvdff #(.WIDTH(1)) dccm_wrbyp_dm_loff(
				.rst_l(rst_l),
				.din(dccm_wr_bypass_d_m_lo),
				.dout(dccm_wr_bypass_d_m_lo_Q),
				.clk(lsu_free_c2_clk)
			);
			rvdff #(.WIDTH(1)) dccm_wrbyp_dm_hiff(
				.rst_l(rst_l),
				.din(dccm_wr_bypass_d_m_hi),
				.dout(dccm_wr_bypass_d_m_hi_Q),
				.clk(lsu_free_c2_clk)
			);
			rvdff #(.WIDTH(32)) store_data_rff(
				.rst_l(rst_l),
				.din(store_data_m[31:0]),
				.dout(store_data_r[31:0]),
				.clk(lsu_store_c1_r_clk)
			);
		end
		else begin : L2U1_Plus1_0
			wire [31:0] store_data_hi_m;
			wire [31:0] store_data_lo_m;
			wire [63:0] store_data_mask;
			assign {store_data_hi_m[31:0], store_data_lo_m[31:0]} = {32'b00000000000000000000000000000000, store_data_m[31:0]} << (8 * lsu_addr_m[1:0]);
			genvar i;
			for (i = 0; i < 4; i = i + 1) begin
				assign store_data_hi_r_in[(8 * i) + 7:8 * i] = (store_byteen_ext_m[i + 4] ? store_data_hi_m[(8 * i) + 7:8 * i] : (lsu_stbuf_commit_any & dccm_wr_bypass_d_m_hi ? stbuf_data_any[(8 * i) + 7:8 * i] : sec_data_hi_m[(8 * i) + 7:8 * i]));
				assign store_data_lo_r_in[(8 * i) + 7:8 * i] = (store_byteen_ext_m[i] ? store_data_lo_m[(8 * i) + 7:8 * i] : (lsu_stbuf_commit_any & dccm_wr_bypass_d_m_lo ? stbuf_data_any[(8 * i) + 7:8 * i] : sec_data_lo_m[(8 * i) + 7:8 * i]));
				assign store_datafn_lo_r[(8 * i) + 7:8 * i] = ((lsu_stbuf_commit_any & dccm_wr_bypass_d_r_lo) & ~store_byteen_ext_r[i] ? stbuf_data_any[(8 * i) + 7:8 * i] : store_data_lo_r[(8 * i) + 7:8 * i]);
				assign store_datafn_hi_r[(8 * i) + 7:8 * i] = ((lsu_stbuf_commit_any & dccm_wr_bypass_d_r_hi) & ~store_byteen_ext_r[i + 4] ? stbuf_data_any[(8 * i) + 7:8 * i] : store_data_hi_r[(8 * i) + 7:8 * i]);
			end
			for (i = 0; i < 4; i = i + 1) assign store_data_mask[(8 * i) + 7:8 * i] = {8 {store_byteen_r[i]}};
			function automatic [31:0] sv2v_cast_32;
				input reg [31:0] inp;
				sv2v_cast_32 = inp;
			endfunction
			assign store_data_r[31:0] = sv2v_cast_32({store_data_hi_r[31:0], store_data_lo_r[31:0]} >> (8 * lsu_addr_r[1:0])) & store_data_mask[31:0];
			rvdffe #(.WIDTH(pt[1382-:10])) store_data_hi_rff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(store_data_hi_r_in[pt[1382-:10] - 1:0]),
				.dout(store_data_hi_r[pt[1382-:10] - 1:0]),
				.en(((ldst_dual_m & lsu_pkt_m[0]) & lsu_pkt_m[6]) | clk_override),
				.clk(clk)
			);
			rvdff #(.WIDTH(pt[1382-:10])) store_data_lo_rff(
				.rst_l(rst_l),
				.din(store_data_lo_r_in[pt[1382-:10] - 1:0]),
				.dout(store_data_lo_r[pt[1382-:10] - 1:0]),
				.clk(lsu_store_c1_r_clk)
			);
		end
	endgenerate
	assign dccm_rdata_lo_m[pt[1382-:10] - 1:0] = dccm_rd_data_lo[pt[1382-:10] - 1:0];
	assign dccm_rdata_hi_m[pt[1382-:10] - 1:0] = dccm_rd_data_hi[pt[1382-:10] - 1:0];
	assign dccm_data_ecc_lo_m[pt[1372-:7] - 1:0] = dccm_rd_data_lo[pt[1360-:10] - 1:pt[1382-:10]];
	assign dccm_data_ecc_hi_m[pt[1372-:7] - 1:0] = dccm_rd_data_hi[pt[1360-:10] - 1:pt[1382-:10]];
	assign picm_wren = (((lsu_pkt_r[0] & lsu_pkt_r[6]) & addr_in_pic_r) & lsu_commit_r) | dma_pic_wen;
	assign picm_rden = (lsu_pkt_d[0] & lsu_pkt_d[7]) & addr_in_pic_d;
	assign picm_mken = (lsu_pkt_d[0] & lsu_pkt_d[6]) & addr_in_pic_d;
	assign picm_rdaddr[31:0] = pt[130-:36] | {{32 - pt[94-:9] {1'b0}}, lsu_addr_d[pt[94-:9] - 1:0]};
	assign picm_wraddr[31:0] = pt[130-:36] | {{32 - pt[94-:9] {1'b0}}, (dma_pic_wen ? dma_mem_addr[pt[94-:9] - 1:0] : lsu_addr_r[pt[94-:9] - 1:0])};
	assign picm_wr_data[31:0] = (dma_pic_wen ? dma_mem_wdata[31:0] : store_datafn_lo_r[31:0]);
	assign picm_mask_data_m[31:0] = picm_rd_data_m[31:0];
	assign picm_rd_data_m[63:0] = {picm_rd_data[31:0], picm_rd_data[31:0]};
	generate
		if (pt[1365-:5] == 1) begin : Gen_dccm_enable
			rvdff #(.WIDTH(1)) dccm_rden_mff(
				.rst_l(rst_l),
				.din(lsu_dccm_rden_d),
				.dout(lsu_dccm_rden_m),
				.clk(lsu_c2_m_clk)
			);
			rvdff #(.WIDTH(1)) dccm_rden_rff(
				.rst_l(rst_l),
				.din(lsu_dccm_rden_m),
				.dout(lsu_dccm_rden_r),
				.clk(lsu_c2_r_clk)
			);
			rvdff #(.WIDTH(1)) ld_double_ecc_error_rff(
				.rst_l(rst_l),
				.din(lsu_double_ecc_error_r),
				.dout(lsu_double_ecc_error_r_ff),
				.clk(lsu_free_c2_clk)
			);
			rvdff #(.WIDTH(1)) ld_single_ecc_error_hi_rff(
				.rst_l(rst_l),
				.din(ld_single_ecc_error_hi_r_ns),
				.dout(ld_single_ecc_error_hi_r_ff),
				.clk(lsu_free_c2_clk)
			);
			rvdff #(.WIDTH(1)) ld_single_ecc_error_lo_rff(
				.rst_l(rst_l),
				.din(ld_single_ecc_error_lo_r_ns),
				.dout(ld_single_ecc_error_lo_r_ff),
				.clk(lsu_free_c2_clk)
			);
			rvdffe #(.WIDTH(pt[1398-:9])) ld_sec_addr_hi_rff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(end_addr_r[pt[1398-:9] - 1:0]),
				.dout(ld_sec_addr_hi_r_ff[pt[1398-:9] - 1:0]),
				.en(ld_single_ecc_error_r | clk_override),
				.clk(clk)
			);
			rvdffe #(.WIDTH(pt[1398-:9])) ld_sec_addr_lo_rff(
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(lsu_addr_r[pt[1398-:9] - 1:0]),
				.dout(ld_sec_addr_lo_r_ff[pt[1398-:9] - 1:0]),
				.en(ld_single_ecc_error_r | clk_override),
				.clk(clk)
			);
		end
		else begin : Gen_dccm_disable
			assign lsu_dccm_rden_m = 1'b0;
			assign lsu_dccm_rden_r = 1'b0;
			assign lsu_double_ecc_error_r_ff = 1'b0;
			assign ld_single_ecc_error_hi_r_ff = 1'b0;
			assign ld_single_ecc_error_lo_r_ff = 1'b0;
			assign ld_sec_addr_hi_r_ff[pt[1398-:9] - 1:0] = {pt[1398-:9] {1'sb0}};
			assign ld_sec_addr_lo_r_ff[pt[1398-:9] - 1:0] = {pt[1398-:9] {1'sb0}};
		end
	endgenerate
endmodule
module eb1_lsu_dccm_mem (
`ifdef USE_POWER_PINS	
	VPWR,
	VGND,
`endif
	clk,
	active_clk,
	rst_l,
	clk_override,
	dccm_wren,
	dccm_rden,
	dccm_wr_addr_lo,
	dccm_wr_addr_hi,
	dccm_rd_addr_lo,
	dccm_rd_addr_hi,
	dccm_wr_data_lo,
	dccm_wr_data_hi,
	dccm_ext_in_pkt,
	dccm_rd_data_lo,
	dccm_rd_data_hi,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
`ifdef USE_POWER_PINS
	inout wire VPWR;
	inout wire VGND;
`endif
	input wire clk;
	input wire active_clk;
	input wire rst_l;
	input wire clk_override;
	input wire dccm_wren;
	input wire dccm_rden;
	input wire [pt[1398-:9] - 1:0] dccm_wr_addr_lo;
	input wire [pt[1398-:9] - 1:0] dccm_wr_addr_hi;
	input wire [pt[1398-:9] - 1:0] dccm_rd_addr_lo;
	input wire [pt[1398-:9] - 1:0] dccm_rd_addr_hi;
	input wire [pt[1360-:10] - 1:0] dccm_wr_data_lo;
	input wire [pt[1360-:10] - 1:0] dccm_wr_data_hi;
	input wire [(pt[1342-:9] * 12) - 1:0] dccm_ext_in_pkt;
	output wire [pt[1360-:10] - 1:0] dccm_rd_data_lo;
	output wire [pt[1360-:10] - 1:0] dccm_rd_data_hi;
	input wire scan_mode;
	localparam DCCM_WIDTH_BITS = $clog2(pt[1389-:7]);
	localparam DCCM_INDEX_BITS = (pt[1398-:9] - pt[1405-:7]) - pt[1275-:6];
	localparam DCCM_INDEX_DEPTH = (pt[1289-:14] * 1024) / (pt[1389-:7] * pt[1342-:9]);
	wire [pt[1342-:9] - 1:0] wren_bank;
	wire [pt[1342-:9] - 1:0] rden_bank;
	wire [((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? (pt[1342-:9] * (((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1)) + (pt[1405-:7] + 1) : (pt[1342-:9] * (((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)) + (pt[1398-:9] - 2)):((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1)] addr_bank;
	wire [pt[1398-:9] - 1:pt[1405-:7] + DCCM_WIDTH_BITS] rd_addr_even;
	wire [pt[1398-:9] - 1:pt[1405-:7] + DCCM_WIDTH_BITS] rd_addr_odd;
	wire rd_unaligned;
	wire wr_unaligned;
	wire [(pt[1342-:9] * pt[1360-:10]) - 1:0] dccm_bank_dout;
	wire [pt[1360-:10] - 1:0] wrdata;
	wire [(pt[1342-:9] * pt[1360-:10]) - 1:0] wr_data_bank;
	wire [(DCCM_WIDTH_BITS + pt[1405-:7]) - 1:DCCM_WIDTH_BITS] dccm_rd_addr_lo_q;
	wire [(DCCM_WIDTH_BITS + pt[1405-:7]) - 1:DCCM_WIDTH_BITS] dccm_rd_addr_hi_q;
	wire [pt[1342-:9] - 1:0] dccm_clken;
	assign rd_unaligned = dccm_rd_addr_lo[DCCM_WIDTH_BITS+:pt[1405-:7]] != dccm_rd_addr_hi[DCCM_WIDTH_BITS+:pt[1405-:7]];
	assign wr_unaligned = dccm_wr_addr_lo[DCCM_WIDTH_BITS+:pt[1405-:7]] != dccm_wr_addr_hi[DCCM_WIDTH_BITS+:pt[1405-:7]];
	assign dccm_rd_data_lo[pt[1360-:10] - 1:0] = dccm_bank_dout[(dccm_rd_addr_lo_q[pt[1275-:6]+:pt[1405-:7]] * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]];
	assign dccm_rd_data_hi[pt[1360-:10] - 1:0] = dccm_bank_dout[(dccm_rd_addr_hi_q[DCCM_WIDTH_BITS+:pt[1405-:7]] * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]];
	generate
		genvar i;
		for (i = 0; i < pt[1342-:9]; i = i + 1) begin : mem_bank
			assign wren_bank[i] = dccm_wren & ((dccm_wr_addr_hi[2+:pt[1405-:7]] == i) | (dccm_wr_addr_lo[2+:pt[1405-:7]] == i));
			assign rden_bank[i] = dccm_rden & ((dccm_rd_addr_hi[2+:pt[1405-:7]] == i) | (dccm_rd_addr_lo[2+:pt[1405-:7]] == i));
			assign addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)) + ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + DCCM_WIDTH_BITS : (pt[1405-:7] + 2) - ((pt[1405-:7] + DCCM_WIDTH_BITS) - (pt[1398-:9] - 1))) : (((i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)) + ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + DCCM_WIDTH_BITS : (pt[1405-:7] + 2) - ((pt[1405-:7] + DCCM_WIDTH_BITS) - (pt[1398-:9] - 1)))) - DCCM_INDEX_BITS) + 1)+:DCCM_INDEX_BITS] = (wren_bank[i] ? ((dccm_wr_addr_hi[2+:pt[1405-:7]] == i) & wr_unaligned ? dccm_wr_addr_hi[pt[1405-:7] + DCCM_WIDTH_BITS+:DCCM_INDEX_BITS] : dccm_wr_addr_lo[pt[1405-:7] + DCCM_WIDTH_BITS+:DCCM_INDEX_BITS]) : ((dccm_rd_addr_hi[2+:pt[1405-:7]] == i) & rd_unaligned ? dccm_rd_addr_hi[pt[1405-:7] + DCCM_WIDTH_BITS+:DCCM_INDEX_BITS] : dccm_rd_addr_lo[pt[1405-:7] + DCCM_WIDTH_BITS+:DCCM_INDEX_BITS]));
			assign wr_data_bank[i * pt[1360-:10]+:pt[1360-:10]] = ((dccm_wr_addr_hi[2+:pt[1405-:7]] == i) & wr_unaligned ? dccm_wr_data_hi[pt[1360-:10] - 1:0] : dccm_wr_data_lo[pt[1360-:10] - 1:0]);
			assign dccm_clken[i] = (wren_bank[i] | rden_bank[i]) | clk_override;
			if (DCCM_INDEX_DEPTH == 32768) begin : dccm
				ram_32768x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 16384) begin : dccm
				ram_16384x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 8192) begin : dccm
				ram_8192x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 4096) begin : dccm
				ram_4096x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 3072) begin : dccm
				ram_3072x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 2048) begin : dccm
				ram_2048x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 1024) begin : dccm
				sky130_sram_1kbyte_1rw1r_32x256_8 sram(
					`ifdef USE_POWER_PINS
					.vccd1(VPWR),
					.vssd1(VGND),
					`endif
					.clk0(clk),
					.csb0(~dccm_clken[i]),
					.web0(~wren_bank[i]),
					.wmask0(4'hf),
					.addr0(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.din0(wr_data_bank[i * pt[1360-:10]+:pt[1360-:10]]),
					.dout0(dccm_bank_dout[i * pt[1360-:10]+:pt[1360-:10]]),
					.clk1(clk),
					.csb1(1'b1),
					.addr1(8'h00),
					.dout1()
				);
			end
			else if (DCCM_INDEX_DEPTH == 512) begin : dccm
				ram_512x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
			else if (DCCM_INDEX_DEPTH == 256) begin : dccm
				sky130_sram_1kbyte_1rw1r_32x256_8 sram(
					`ifdef USE_POWER_PINS
					.vccd1(VPWR),
					.vssd1(VGND),
					`endif
					.clk0(clk),
					.csb0(~dccm_clken[i]),
					.web0(~wren_bank[i]),
					.wmask0(4'hf),
					.addr0(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.din0(wr_data_bank[(i * pt[1360-:10]) + 31-:32]),
					.dout0(dccm_bank_dout[(i * pt[1360-:10]) + 31-:32]),
					.clk1(clk),
					.csb1(1'b1),
					.addr1(8'h00),
					.dout1()
				);
			end
			else if (DCCM_INDEX_DEPTH == 128) begin : dccm
				ram_128x39 dccm_bank(
					.ME(dccm_clken[i]),
					.CLK(clk),
					.WE(wren_bank[i]),
					.ADR(addr_bank[((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? pt[1405-:7] + 2 : pt[1398-:9] - 1) + (i * ((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1))+:((pt[1398-:9] - 1) >= (pt[1405-:7] + 2) ? ((pt[1398-:9] - 1) - (pt[1405-:7] + 2)) + 1 : ((pt[1405-:7] + 2) - (pt[1398-:9] - 1)) + 1)]),
					.D(wr_data_bank[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.Q(dccm_bank_dout[(i * pt[1360-:10]) + (pt[1360-:10] - 1)-:pt[1360-:10]]),
					.ROP(),
					.TEST1(dccm_ext_in_pkt[(i * 12) + 11]),
					.RME(dccm_ext_in_pkt[(i * 12) + 10]),
					.RM(dccm_ext_in_pkt[(i * 12) + 9-:4]),
					.LS(dccm_ext_in_pkt[(i * 12) + 5]),
					.DS(dccm_ext_in_pkt[(i * 12) + 4]),
					.SD(dccm_ext_in_pkt[(i * 12) + 3]),
					.TEST_RNM(dccm_ext_in_pkt[(i * 12) + 2]),
					.BC1(dccm_ext_in_pkt[(i * 12) + 1]),
					.BC2(dccm_ext_in_pkt[i * 12]),
					.*
				);
			end
		end
	endgenerate
	rvdff #(.WIDTH(pt[1405-:7])) rd_addr_lo_ff(
		.rst_l(rst_l),
		.din(dccm_rd_addr_lo[DCCM_WIDTH_BITS+:pt[1405-:7]]),
		.dout(dccm_rd_addr_lo_q[DCCM_WIDTH_BITS+:pt[1405-:7]]),
		.clk(active_clk)
	);
	rvdff #(.WIDTH(pt[1405-:7])) rd_addr_hi_ff(
		.rst_l(rst_l),
		.din(dccm_rd_addr_hi[DCCM_WIDTH_BITS+:pt[1405-:7]]),
		.dout(dccm_rd_addr_hi_q[DCCM_WIDTH_BITS+:pt[1405-:7]]),
		.clk(active_clk)
	);
endmodule
module eb1_lsu_ecc (
	clk,
	lsu_c2_r_clk,
	clk_override,
	rst_l,
	scan_mode,
	lsu_pkt_m,
	lsu_pkt_r,
	stbuf_data_any,
	dec_tlu_core_ecc_disable,
	lsu_dccm_rden_r,
	addr_in_dccm_r,
	lsu_addr_r,
	end_addr_r,
	dccm_rdata_hi_r,
	dccm_rdata_lo_r,
	dccm_data_ecc_hi_r,
	dccm_data_ecc_lo_r,
	sec_data_hi_r,
	sec_data_lo_r,
	sec_data_hi_r_ff,
	sec_data_lo_r_ff,
	ld_single_ecc_error_r,
	ld_single_ecc_error_r_ff,
	lsu_dccm_rden_m,
	addr_in_dccm_m,
	lsu_addr_m,
	end_addr_m,
	dccm_rdata_hi_m,
	dccm_rdata_lo_m,
	dccm_data_ecc_hi_m,
	dccm_data_ecc_lo_m,
	sec_data_hi_m,
	sec_data_lo_m,
	dma_dccm_wen,
	dma_dccm_wdata_lo,
	dma_dccm_wdata_hi,
	dma_dccm_wdata_ecc_hi,
	dma_dccm_wdata_ecc_lo,
	stbuf_ecc_any,
	sec_data_ecc_hi_r_ff,
	sec_data_ecc_lo_r_ff,
	single_ecc_error_hi_r,
	single_ecc_error_lo_r,
	lsu_single_ecc_error_r,
	lsu_double_ecc_error_r,
	lsu_single_ecc_error_m,
	lsu_double_ecc_error_m
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire lsu_c2_r_clk;
	input wire clk_override;
	input wire rst_l;
	input wire scan_mode;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_r;
	input wire [pt[1382-:10] - 1:0] stbuf_data_any;
	input wire dec_tlu_core_ecc_disable;
	input wire lsu_dccm_rden_r;
	input wire addr_in_dccm_r;
	input wire [pt[1398-:9] - 1:0] lsu_addr_r;
	input wire [pt[1398-:9] - 1:0] end_addr_r;
	input wire [pt[1382-:10] - 1:0] dccm_rdata_hi_r;
	input wire [pt[1382-:10] - 1:0] dccm_rdata_lo_r;
	input wire [pt[1372-:7] - 1:0] dccm_data_ecc_hi_r;
	input wire [pt[1372-:7] - 1:0] dccm_data_ecc_lo_r;
	output wire [pt[1382-:10] - 1:0] sec_data_hi_r;
	output wire [pt[1382-:10] - 1:0] sec_data_lo_r;
	output wire [pt[1382-:10] - 1:0] sec_data_hi_r_ff;
	output wire [pt[1382-:10] - 1:0] sec_data_lo_r_ff;
	input wire ld_single_ecc_error_r;
	input wire ld_single_ecc_error_r_ff;
	input wire lsu_dccm_rden_m;
	input wire addr_in_dccm_m;
	input wire [pt[1398-:9] - 1:0] lsu_addr_m;
	input wire [pt[1398-:9] - 1:0] end_addr_m;
	input wire [pt[1382-:10] - 1:0] dccm_rdata_hi_m;
	input wire [pt[1382-:10] - 1:0] dccm_rdata_lo_m;
	input wire [pt[1372-:7] - 1:0] dccm_data_ecc_hi_m;
	input wire [pt[1372-:7] - 1:0] dccm_data_ecc_lo_m;
	output wire [pt[1382-:10] - 1:0] sec_data_hi_m;
	output wire [pt[1382-:10] - 1:0] sec_data_lo_m;
	input wire dma_dccm_wen;
	input wire [31:0] dma_dccm_wdata_lo;
	input wire [31:0] dma_dccm_wdata_hi;
	output wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_hi;
	output wire [pt[1372-:7] - 1:0] dma_dccm_wdata_ecc_lo;
	output wire [pt[1372-:7] - 1:0] stbuf_ecc_any;
	output wire [pt[1372-:7] - 1:0] sec_data_ecc_hi_r_ff;
	output wire [pt[1372-:7] - 1:0] sec_data_ecc_lo_r_ff;
	output wire single_ecc_error_hi_r;
	output wire single_ecc_error_lo_r;
	output wire lsu_single_ecc_error_r;
	output wire lsu_double_ecc_error_r;
	output wire lsu_single_ecc_error_m;
	output wire lsu_double_ecc_error_m;
	wire is_ldst_r;
	wire is_ldst_hi_any;
	wire is_ldst_lo_any;
	wire [pt[1382-:10] - 1:0] dccm_wdata_hi_any;
	wire [pt[1382-:10] - 1:0] dccm_wdata_lo_any;
	wire [pt[1372-:7] - 1:0] dccm_wdata_ecc_hi_any;
	wire [pt[1372-:7] - 1:0] dccm_wdata_ecc_lo_any;
	wire [pt[1382-:10] - 1:0] dccm_rdata_hi_any;
	wire [pt[1382-:10] - 1:0] dccm_rdata_lo_any;
	wire [pt[1372-:7] - 1:0] dccm_data_ecc_hi_any;
	wire [pt[1372-:7] - 1:0] dccm_data_ecc_lo_any;
	wire [pt[1382-:10] - 1:0] sec_data_hi_any;
	wire [pt[1382-:10] - 1:0] sec_data_lo_any;
	wire single_ecc_error_hi_any;
	wire single_ecc_error_lo_any;
	wire double_ecc_error_hi_any;
	wire double_ecc_error_lo_any;
	wire double_ecc_error_hi_m;
	wire double_ecc_error_lo_m;
	wire double_ecc_error_hi_r;
	wire double_ecc_error_lo_r;
	wire [6:0] ecc_out_hi_nc;
	wire [6:0] ecc_out_lo_nc;
	generate
		if (pt[202-:5] == 1) begin : L2U_Plus1_1
			wire ldst_dual_m;
			wire ldst_dual_r;
			wire is_ldst_m;
			wire is_ldst_hi_r;
			wire is_ldst_lo_r;
			assign ldst_dual_r = lsu_addr_r[2] != end_addr_r[2];
			assign is_ldst_r = ((lsu_pkt_r[0] & (lsu_pkt_r[7] | lsu_pkt_r[6])) & addr_in_dccm_r) & lsu_dccm_rden_r;
			assign is_ldst_lo_r = is_ldst_r & ~dec_tlu_core_ecc_disable;
			assign is_ldst_hi_r = (is_ldst_r & ldst_dual_r) & ~dec_tlu_core_ecc_disable;
			assign is_ldst_hi_any = is_ldst_hi_r;
			assign dccm_rdata_hi_any[pt[1382-:10] - 1:0] = dccm_rdata_hi_r[pt[1382-:10] - 1:0];
			assign dccm_data_ecc_hi_any[pt[1372-:7] - 1:0] = dccm_data_ecc_hi_r[pt[1372-:7] - 1:0];
			assign is_ldst_lo_any = is_ldst_lo_r;
			assign dccm_rdata_lo_any[pt[1382-:10] - 1:0] = dccm_rdata_lo_r[pt[1382-:10] - 1:0];
			assign dccm_data_ecc_lo_any[pt[1372-:7] - 1:0] = dccm_data_ecc_lo_r[pt[1372-:7] - 1:0];
			assign sec_data_hi_r[pt[1382-:10] - 1:0] = sec_data_hi_any[pt[1382-:10] - 1:0];
			assign single_ecc_error_hi_r = single_ecc_error_hi_any;
			assign double_ecc_error_hi_r = double_ecc_error_hi_any;
			assign sec_data_lo_r[pt[1382-:10] - 1:0] = sec_data_lo_any[pt[1382-:10] - 1:0];
			assign single_ecc_error_lo_r = single_ecc_error_lo_any;
			assign double_ecc_error_lo_r = double_ecc_error_lo_any;
			assign lsu_single_ecc_error_r = single_ecc_error_hi_r | single_ecc_error_lo_r;
			assign lsu_double_ecc_error_r = double_ecc_error_hi_r | double_ecc_error_lo_r;
		end
		else begin : L2U_Plus1_0
			wire ldst_dual_m;
			wire is_ldst_m;
			wire is_ldst_hi_m;
			wire is_ldst_lo_m;
			assign ldst_dual_m = lsu_addr_m[2] != end_addr_m[2];
			assign is_ldst_m = ((lsu_pkt_m[0] & (lsu_pkt_m[7] | lsu_pkt_m[6])) & addr_in_dccm_m) & lsu_dccm_rden_m;
			assign is_ldst_lo_m = is_ldst_m & ~dec_tlu_core_ecc_disable;
			assign is_ldst_hi_m = (is_ldst_m & (ldst_dual_m | lsu_pkt_m[4])) & ~dec_tlu_core_ecc_disable;
			assign is_ldst_hi_any = is_ldst_hi_m;
			assign dccm_rdata_hi_any[pt[1382-:10] - 1:0] = dccm_rdata_hi_m[pt[1382-:10] - 1:0];
			assign dccm_data_ecc_hi_any[pt[1372-:7] - 1:0] = dccm_data_ecc_hi_m[pt[1372-:7] - 1:0];
			assign is_ldst_lo_any = is_ldst_lo_m;
			assign dccm_rdata_lo_any[pt[1382-:10] - 1:0] = dccm_rdata_lo_m[pt[1382-:10] - 1:0];
			assign dccm_data_ecc_lo_any[pt[1372-:7] - 1:0] = dccm_data_ecc_lo_m[pt[1372-:7] - 1:0];
			assign sec_data_hi_m[pt[1382-:10] - 1:0] = sec_data_hi_any[pt[1382-:10] - 1:0];
			assign double_ecc_error_hi_m = double_ecc_error_hi_any;
			assign sec_data_lo_m[pt[1382-:10] - 1:0] = sec_data_lo_any[pt[1382-:10] - 1:0];
			assign double_ecc_error_lo_m = double_ecc_error_lo_any;
			assign lsu_single_ecc_error_m = single_ecc_error_hi_any | single_ecc_error_lo_any;
			assign lsu_double_ecc_error_m = double_ecc_error_hi_m | double_ecc_error_lo_m;
			rvdff #(.WIDTH(1)) lsu_single_ecc_err_r(
				.din(lsu_single_ecc_error_m),
				.dout(lsu_single_ecc_error_r),
				.clk(lsu_c2_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) lsu_double_ecc_err_r(
				.din(lsu_double_ecc_error_m),
				.dout(lsu_double_ecc_error_r),
				.clk(lsu_c2_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) ldst_sec_lo_rff(
				.din(single_ecc_error_lo_any),
				.dout(single_ecc_error_lo_r),
				.clk(lsu_c2_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) ldst_sec_hi_rff(
				.din(single_ecc_error_hi_any),
				.dout(single_ecc_error_hi_r),
				.clk(lsu_c2_r_clk),
				.rst_l(rst_l)
			);
			rvdffe #(.WIDTH(pt[1382-:10])) sec_data_hi_rff(
				.din(sec_data_hi_m[pt[1382-:10] - 1:0]),
				.dout(sec_data_hi_r[pt[1382-:10] - 1:0]),
				.en(lsu_single_ecc_error_m | clk_override),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
			rvdffe #(.WIDTH(pt[1382-:10])) sec_data_lo_rff(
				.din(sec_data_lo_m[pt[1382-:10] - 1:0]),
				.dout(sec_data_lo_r[pt[1382-:10] - 1:0]),
				.en(lsu_single_ecc_error_m | clk_override),
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode)
			);
		end
	endgenerate
	assign dccm_wdata_lo_any[pt[1382-:10] - 1:0] = (ld_single_ecc_error_r_ff ? sec_data_lo_r_ff[pt[1382-:10] - 1:0] : (dma_dccm_wen ? dma_dccm_wdata_lo[pt[1382-:10] - 1:0] : stbuf_data_any[pt[1382-:10] - 1:0]));
	assign dccm_wdata_hi_any[pt[1382-:10] - 1:0] = (ld_single_ecc_error_r_ff ? sec_data_hi_r_ff[pt[1382-:10] - 1:0] : (dma_dccm_wen ? dma_dccm_wdata_hi[pt[1382-:10] - 1:0] : 32'h00000000));
	assign sec_data_ecc_hi_r_ff[pt[1372-:7] - 1:0] = dccm_wdata_ecc_hi_any[pt[1372-:7] - 1:0];
	assign sec_data_ecc_lo_r_ff[pt[1372-:7] - 1:0] = dccm_wdata_ecc_lo_any[pt[1372-:7] - 1:0];
	assign stbuf_ecc_any[pt[1372-:7] - 1:0] = dccm_wdata_ecc_lo_any[pt[1372-:7] - 1:0];
	assign dma_dccm_wdata_ecc_hi[pt[1372-:7] - 1:0] = dccm_wdata_ecc_hi_any[pt[1372-:7] - 1:0];
	assign dma_dccm_wdata_ecc_lo[pt[1372-:7] - 1:0] = dccm_wdata_ecc_lo_any[pt[1372-:7] - 1:0];
	generate
		if (pt[1365-:5] == 1) begin : Gen_dccm_enable
			rvecc_decode lsu_ecc_decode_hi(
				.en(is_ldst_hi_any),
				.sed_ded(1'b0),
				.din(dccm_rdata_hi_any[pt[1382-:10] - 1:0]),
				.ecc_in(dccm_data_ecc_hi_any[pt[1372-:7] - 1:0]),
				.dout(sec_data_hi_any[pt[1382-:10] - 1:0]),
				.ecc_out(ecc_out_hi_nc[6:0]),
				.single_ecc_error(single_ecc_error_hi_any),
				.double_ecc_error(double_ecc_error_hi_any)
			);
			rvecc_decode lsu_ecc_decode_lo(
				.en(is_ldst_lo_any),
				.sed_ded(1'b0),
				.din(dccm_rdata_lo_any[pt[1382-:10] - 1:0]),
				.ecc_in(dccm_data_ecc_lo_any[pt[1372-:7] - 1:0]),
				.dout(sec_data_lo_any[pt[1382-:10] - 1:0]),
				.ecc_out(ecc_out_lo_nc[6:0]),
				.single_ecc_error(single_ecc_error_lo_any),
				.double_ecc_error(double_ecc_error_lo_any)
			);
			rvecc_encode lsu_ecc_encode_hi(
				.din(dccm_wdata_hi_any[pt[1382-:10] - 1:0]),
				.ecc_out(dccm_wdata_ecc_hi_any[pt[1372-:7] - 1:0])
			);
			rvecc_encode lsu_ecc_encode_lo(
				.din(dccm_wdata_lo_any[pt[1382-:10] - 1:0]),
				.ecc_out(dccm_wdata_ecc_lo_any[pt[1372-:7] - 1:0])
			);
		end
		else begin : Gen_dccm_disable
			assign sec_data_hi_any[pt[1382-:10] - 1:0] = {pt[1382-:10] {1'sb0}};
			assign sec_data_lo_any[pt[1382-:10] - 1:0] = {pt[1382-:10] {1'sb0}};
			assign single_ecc_error_hi_any = 1'b0;
			assign double_ecc_error_hi_any = 1'b0;
			assign single_ecc_error_lo_any = 1'b0;
			assign double_ecc_error_lo_any = 1'b0;
		end
	endgenerate
	rvdffe #(.WIDTH(pt[1382-:10])) sec_data_hi_rplus1ff(
		.din(sec_data_hi_r[pt[1382-:10] - 1:0]),
		.dout(sec_data_hi_r_ff[pt[1382-:10] - 1:0]),
		.en(ld_single_ecc_error_r | clk_override),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
	rvdffe #(.WIDTH(pt[1382-:10])) sec_data_lo_rplus1ff(
		.din(sec_data_lo_r[pt[1382-:10] - 1:0]),
		.dout(sec_data_lo_r_ff[pt[1382-:10] - 1:0]),
		.en(ld_single_ecc_error_r | clk_override),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode)
	);
endmodule
module eb1_lsu_lsc_ctl (
	rst_l,
	clk_override,
	clk,
	lsu_c1_m_clk,
	lsu_c1_r_clk,
	lsu_c2_m_clk,
	lsu_c2_r_clk,
	lsu_store_c1_m_clk,
	lsu_ld_data_r,
	lsu_ld_data_corr_r,
	lsu_single_ecc_error_r,
	lsu_double_ecc_error_r,
	lsu_ld_data_m,
	lsu_single_ecc_error_m,
	lsu_double_ecc_error_m,
	flush_m_up,
	flush_r,
	ldst_dual_d,
	ldst_dual_m,
	ldst_dual_r,
	exu_lsu_rs1_d,
	exu_lsu_rs2_d,
	lsu_p,
	dec_lsu_valid_raw_d,
	dec_lsu_offset_d,
	picm_mask_data_m,
	bus_read_data_m,
	lsu_result_m,
	lsu_result_corr_r,
	lsu_addr_d,
	lsu_addr_m,
	lsu_addr_r,
	end_addr_d,
	end_addr_m,
	end_addr_r,
	store_data_m,
	dec_tlu_mrac_ff,
	lsu_exc_m,
	is_sideeffects_m,
	lsu_commit_r,
	lsu_single_ecc_error_incr,
	lsu_error_pkt_r,
	lsu_fir_addr,
	lsu_fir_error,
	addr_in_dccm_d,
	addr_in_dccm_m,
	addr_in_dccm_r,
	addr_in_pic_d,
	addr_in_pic_m,
	addr_in_pic_r,
	addr_external_m,
	dma_dccm_req,
	dma_mem_addr,
	dma_mem_sz,
	dma_mem_write,
	dma_mem_wdata,
	lsu_pkt_d,
	lsu_pkt_m,
	lsu_pkt_r,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire rst_l;
	input wire clk_override;
	input wire clk;
	input wire lsu_c1_m_clk;
	input wire lsu_c1_r_clk;
	input wire lsu_c2_m_clk;
	input wire lsu_c2_r_clk;
	input wire lsu_store_c1_m_clk;
	input wire [31:0] lsu_ld_data_r;
	input wire [31:0] lsu_ld_data_corr_r;
	input wire lsu_single_ecc_error_r;
	input wire lsu_double_ecc_error_r;
	input wire [31:0] lsu_ld_data_m;
	input wire lsu_single_ecc_error_m;
	input wire lsu_double_ecc_error_m;
	input wire flush_m_up;
	input wire flush_r;
	input wire ldst_dual_d;
	input wire ldst_dual_m;
	input wire ldst_dual_r;
	input wire [31:0] exu_lsu_rs1_d;
	input wire [31:0] exu_lsu_rs2_d;
	input wire [13:0] lsu_p;
	input wire dec_lsu_valid_raw_d;
	input wire [11:0] dec_lsu_offset_d;
	input wire [31:0] picm_mask_data_m;
	input wire [31:0] bus_read_data_m;
	output wire [31:0] lsu_result_m;
	output wire [31:0] lsu_result_corr_r;
	output wire [31:0] lsu_addr_d;
	output wire [31:0] lsu_addr_m;
	output wire [31:0] lsu_addr_r;
	output wire [31:0] end_addr_d;
	output wire [31:0] end_addr_m;
	output wire [31:0] end_addr_r;
	output wire [31:0] store_data_m;
	input wire [31:0] dec_tlu_mrac_ff;
	output wire lsu_exc_m;
	output wire is_sideeffects_m;
	output wire lsu_commit_r;
	output wire lsu_single_ecc_error_incr;
	output wire [39:0] lsu_error_pkt_r;
	output wire [31:1] lsu_fir_addr;
	output wire [1:0] lsu_fir_error;
	output wire addr_in_dccm_d;
	output wire addr_in_dccm_m;
	output wire addr_in_dccm_r;
	output wire addr_in_pic_d;
	output wire addr_in_pic_m;
	output wire addr_in_pic_r;
	output wire addr_external_m;
	input wire dma_dccm_req;
	input wire [31:0] dma_mem_addr;
	input wire [2:0] dma_mem_sz;
	input wire dma_mem_write;
	input wire [63:0] dma_mem_wdata;
	output reg [13:0] lsu_pkt_d;
	output wire [13:0] lsu_pkt_m;
	output wire [13:0] lsu_pkt_r;
	input wire scan_mode;
	wire [31:3] end_addr_pre_m;
	wire [31:3] end_addr_pre_r;
	wire [31:0] full_addr_d;
	wire [31:0] full_end_addr_d;
	wire [31:0] lsu_rs1_d;
	wire [11:0] lsu_offset_d;
	wire [31:0] rs1_d;
	wire [11:0] offset_d;
	wire [12:0] end_addr_offset_d;
	wire [2:0] addr_offset_d;
	wire [63:0] dma_mem_wdata_shifted;
	wire addr_external_d;
	wire addr_external_r;
	wire access_fault_d;
	wire misaligned_fault_d;
	wire access_fault_m;
	wire misaligned_fault_m;
	wire fir_dccm_access_error_d;
	wire fir_nondccm_access_error_d;
	wire fir_dccm_access_error_m;
	wire fir_nondccm_access_error_m;
	wire [3:0] exc_mscause_d;
	wire [3:0] exc_mscause_m;
	wire [31:0] rs1_d_raw;
	wire [31:0] store_data_d;
	wire [31:0] store_data_pre_m;
	wire [31:0] store_data_m_in;
	wire [31:0] bus_read_data_r;
	reg [13:0] dma_pkt_d;
	reg [13:0] lsu_pkt_m_in;
	reg [13:0] lsu_pkt_r_in;
	wire [39:0] lsu_error_pkt_m;
	assign lsu_rs1_d[31:0] = (dec_lsu_valid_raw_d ? exu_lsu_rs1_d[31:0] : dma_mem_addr[31:0]);
	assign lsu_offset_d[11:0] = dec_lsu_offset_d[11:0] & {12 {dec_lsu_valid_raw_d}};
	assign rs1_d_raw[31:0] = lsu_rs1_d[31:0];
	assign offset_d[11:0] = lsu_offset_d[11:0];
	assign rs1_d[31:0] = (lsu_pkt_d[2] ? lsu_result_m[31:0] : rs1_d_raw[31:0]);
	rvlsadder lsadder(
		.rs1(rs1_d[31:0]),
		.offset(offset_d[11:0]),
		.dout(full_addr_d[31:0])
	);
	eb1_lsu_addrcheck #(.pt(pt)) addrcheck(
		.start_addr_d(full_addr_d[31:0]),
		.end_addr_d(full_end_addr_d[31:0]),
		.rs1_region_d(rs1_d[31:28]),
		.lsu_c2_m_clk(lsu_c2_m_clk),
		.rst_l(rst_l),
		.lsu_pkt_d(lsu_pkt_d),
		.dec_tlu_mrac_ff(dec_tlu_mrac_ff),
		.rs1_d(rs1_d),
		.is_sideeffects_m(is_sideeffects_m),
		.addr_in_dccm_d(addr_in_dccm_d),
		.addr_in_pic_d(addr_in_pic_d),
		.addr_external_d(addr_external_d),
		.access_fault_d(access_fault_d),
		.misaligned_fault_d(misaligned_fault_d),
		.exc_mscause_d(exc_mscause_d),
		.fir_dccm_access_error_d(fir_dccm_access_error_d),
		.fir_nondccm_access_error_d(fir_nondccm_access_error_d),
		.scan_mode(scan_mode)
	);
	assign addr_offset_d[2:0] = (({3 {lsu_pkt_d[10]}} & 3'b001) | ({3 {lsu_pkt_d[9]}} & 3'b011)) | ({3 {lsu_pkt_d[8]}} & 3'b111);
	assign end_addr_offset_d[12:0] = {offset_d[11], offset_d[11:0]} + {9'b000000000, addr_offset_d[2:0]};
	assign full_end_addr_d[31:0] = rs1_d[31:0] + {{19 {end_addr_offset_d[12]}}, end_addr_offset_d[12:0]};
	assign end_addr_d[31:0] = full_end_addr_d[31:0];
	assign lsu_exc_m = access_fault_m | misaligned_fault_m;
	assign lsu_single_ecc_error_incr = ((lsu_single_ecc_error_r & ~lsu_double_ecc_error_r) & (lsu_commit_r | lsu_pkt_r[4])) & lsu_pkt_r[0];
	generate
		if (pt[202-:5] == 1) begin : L2U_Plus1_1
			wire access_fault_r;
			wire misaligned_fault_r;
			wire [3:0] exc_mscause_r;
			wire fir_dccm_access_error_r;
			wire fir_nondccm_access_error_r;
			assign lsu_error_pkt_r[0] = ((((access_fault_r | misaligned_fault_r) | lsu_double_ecc_error_r) & lsu_pkt_r[0]) & ~lsu_pkt_r[4]) & ~lsu_pkt_r[13];
			assign lsu_error_pkt_r[1] = (lsu_single_ecc_error_r & ~lsu_error_pkt_r[0]) & ~lsu_pkt_r[4];
			assign lsu_error_pkt_r[39] = lsu_pkt_r[6];
			assign lsu_error_pkt_r[38] = ~misaligned_fault_r;
			assign lsu_error_pkt_r[37:34] = ((lsu_double_ecc_error_r & ~misaligned_fault_r) & ~access_fault_r ? 4'h1 : exc_mscause_r[3:0]);
			assign lsu_error_pkt_r[33:2] = lsu_addr_r[31:0];
			assign lsu_fir_error[1:0] = (fir_nondccm_access_error_r ? 2'b11 : (fir_dccm_access_error_r ? 2'b10 : (lsu_pkt_r[13] & lsu_double_ecc_error_r ? 2'b01 : 2'b00)));
			rvdff #(.WIDTH(1)) access_fault_rff(
				.din(access_fault_m),
				.dout(access_fault_r),
				.clk(lsu_c1_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) misaligned_fault_rff(
				.din(misaligned_fault_m),
				.dout(misaligned_fault_r),
				.clk(lsu_c1_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(4)) exc_mscause_rff(
				.din(exc_mscause_m[3:0]),
				.dout(exc_mscause_r[3:0]),
				.clk(lsu_c1_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) fir_dccm_access_error_mff(
				.din(fir_dccm_access_error_m),
				.dout(fir_dccm_access_error_r),
				.clk(lsu_c1_r_clk),
				.rst_l(rst_l)
			);
			rvdff #(.WIDTH(1)) fir_nondccm_access_error_mff(
				.din(fir_nondccm_access_error_m),
				.dout(fir_nondccm_access_error_r),
				.clk(lsu_c1_r_clk),
				.rst_l(rst_l)
			);
		end
		else begin : L2U_Plus1_0
			wire [1:0] lsu_fir_error_m;
			assign lsu_error_pkt_m[0] = (((((access_fault_m | misaligned_fault_m) | lsu_double_ecc_error_m) & lsu_pkt_m[0]) & ~lsu_pkt_m[4]) & ~lsu_pkt_m[13]) & ~flush_m_up;
			assign lsu_error_pkt_m[1] = (lsu_single_ecc_error_m & ~lsu_error_pkt_m[0]) & ~lsu_pkt_m[4];
			assign lsu_error_pkt_m[39] = lsu_pkt_m[6];
			assign lsu_error_pkt_m[38] = ~misaligned_fault_m;
			assign lsu_error_pkt_m[37:34] = ((lsu_double_ecc_error_m & ~misaligned_fault_m) & ~access_fault_m ? 4'h1 : exc_mscause_m[3:0]);
			assign lsu_error_pkt_m[33:2] = lsu_addr_m[31:0];
			assign lsu_fir_error_m[1:0] = (fir_nondccm_access_error_m ? 2'b11 : (fir_dccm_access_error_m ? 2'b10 : (lsu_pkt_m[13] & lsu_double_ecc_error_m ? 2'b01 : 2'b00)));
			rvdff #(.WIDTH(1)) lsu_exc_valid_rff(
				.rst_l(rst_l),
				.din(lsu_error_pkt_m[0]),
				.dout(lsu_error_pkt_r[0]),
				.clk(lsu_c2_r_clk)
			);
			rvdff #(.WIDTH(1)) lsu_single_ecc_error_rff(
				.rst_l(rst_l),
				.din(lsu_error_pkt_m[1]),
				.dout(lsu_error_pkt_r[1]),
				.clk(lsu_c2_r_clk)
			);
			rvdffe #(.WIDTH(38)) lsu_error_pkt_rff(
				.clk(clk),
				.rst_l(rst_l),
				.scan_mode(scan_mode),
				.din(lsu_error_pkt_m[39:2]),
				.dout(lsu_error_pkt_r[39:2]),
				.en((lsu_error_pkt_m[0] | lsu_error_pkt_m[1]) | clk_override)
			);
			rvdff #(.WIDTH(2)) lsu_fir_error_rff(
				.rst_l(rst_l),
				.din(lsu_fir_error_m[1:0]),
				.dout(lsu_fir_error[1:0]),
				.clk(lsu_c2_r_clk)
			);
		end
	endgenerate
	always @(*) begin
		dma_pkt_d = {14 {1'sb0}};
		dma_pkt_d[0] = dma_dccm_req;
		dma_pkt_d[4] = 1'b1;
		dma_pkt_d[6] = dma_mem_write;
		dma_pkt_d[7] = ~dma_mem_write;
		dma_pkt_d[11] = dma_mem_sz[2:0] == 3'b000;
		dma_pkt_d[10] = dma_mem_sz[2:0] == 3'b001;
		dma_pkt_d[9] = dma_mem_sz[2:0] == 3'b010;
		dma_pkt_d[8] = dma_mem_sz[2:0] == 3'b011;
	end
	always @(*) begin
		lsu_pkt_d = (dec_lsu_valid_raw_d ? lsu_p : dma_pkt_d);
		lsu_pkt_m_in = lsu_pkt_d;
		lsu_pkt_r_in = lsu_pkt_m;
		lsu_pkt_d[0] = (lsu_p[0] & ~(flush_m_up & ~lsu_p[13])) | dma_dccm_req;
		lsu_pkt_m_in[0] = lsu_pkt_d[0] & ~(flush_m_up & ~lsu_pkt_d[4]);
		lsu_pkt_r_in[0] = lsu_pkt_m[0] & ~(flush_m_up & ~lsu_pkt_m[4]);
	end
	rvdff #(.WIDTH(1)) lsu_pkt_vldmff(
		.rst_l(rst_l),
		.din(lsu_pkt_m_in[0]),
		.dout(lsu_pkt_m[0]),
		.clk(lsu_c2_m_clk)
	);
	rvdff #(.WIDTH(1)) lsu_pkt_vldrff(
		.rst_l(rst_l),
		.din(lsu_pkt_r_in[0]),
		.dout(lsu_pkt_r[0]),
		.clk(lsu_c2_r_clk)
	);
	rvdff #(.WIDTH(13)) lsu_pkt_mff(
		.rst_l(rst_l),
		.din(lsu_pkt_m_in[13:1]),
		.dout(lsu_pkt_m[13:1]),
		.clk(lsu_c1_m_clk)
	);
	rvdff #(.WIDTH(13)) lsu_pkt_rff(
		.rst_l(rst_l),
		.din(lsu_pkt_r_in[13:1]),
		.dout(lsu_pkt_r[13:1]),
		.clk(lsu_c1_r_clk)
	);
	generate
		if (pt[202-:5] == 1) begin : L2U1_Plus1_1
			wire [31:0] lsu_ld_datafn_r;
			wire [31:0] lsu_ld_datafn_corr_r;
			assign lsu_ld_datafn_r[31:0] = (addr_external_r ? bus_read_data_r[31:0] : lsu_ld_data_r[31:0]);
			assign lsu_ld_datafn_corr_r[31:0] = (addr_external_r ? bus_read_data_r[31:0] : lsu_ld_data_corr_r[31:0]);
			assign lsu_result_m[31:0] = (((({32 {lsu_pkt_r[5] & lsu_pkt_r[11]}} & {24'b000000000000000000000000, lsu_ld_datafn_r[7:0]}) | ({32 {lsu_pkt_r[5] & lsu_pkt_r[10]}} & {16'b0000000000000000, lsu_ld_datafn_r[15:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[11]}} & {{24 {lsu_ld_datafn_r[7]}}, lsu_ld_datafn_r[7:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[10]}} & {{16 {lsu_ld_datafn_r[15]}}, lsu_ld_datafn_r[15:0]})) | ({32 {lsu_pkt_r[9]}} & lsu_ld_datafn_r[31:0]);
			assign lsu_result_corr_r[31:0] = (((({32 {lsu_pkt_r[5] & lsu_pkt_r[11]}} & {24'b000000000000000000000000, lsu_ld_datafn_corr_r[7:0]}) | ({32 {lsu_pkt_r[5] & lsu_pkt_r[10]}} & {16'b0000000000000000, lsu_ld_datafn_corr_r[15:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[11]}} & {{24 {lsu_ld_datafn_corr_r[7]}}, lsu_ld_datafn_corr_r[7:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[10]}} & {{16 {lsu_ld_datafn_corr_r[15]}}, lsu_ld_datafn_corr_r[15:0]})) | ({32 {lsu_pkt_r[9]}} & lsu_ld_datafn_corr_r[31:0]);
		end
		else begin : L2U1_Plus1_0
			wire [31:0] lsu_ld_datafn_m;
			wire [31:0] lsu_ld_datafn_corr_r;
			assign lsu_ld_datafn_m[31:0] = (addr_external_m ? bus_read_data_m[31:0] : lsu_ld_data_m[31:0]);
			assign lsu_ld_datafn_corr_r[31:0] = (addr_external_r ? bus_read_data_r[31:0] : lsu_ld_data_corr_r[31:0]);
			assign lsu_result_m[31:0] = (((({32 {lsu_pkt_m[5] & lsu_pkt_m[11]}} & {24'b000000000000000000000000, lsu_ld_datafn_m[7:0]}) | ({32 {lsu_pkt_m[5] & lsu_pkt_m[10]}} & {16'b0000000000000000, lsu_ld_datafn_m[15:0]})) | ({32 {~lsu_pkt_m[5] & lsu_pkt_m[11]}} & {{24 {lsu_ld_datafn_m[7]}}, lsu_ld_datafn_m[7:0]})) | ({32 {~lsu_pkt_m[5] & lsu_pkt_m[10]}} & {{16 {lsu_ld_datafn_m[15]}}, lsu_ld_datafn_m[15:0]})) | ({32 {lsu_pkt_m[9]}} & lsu_ld_datafn_m[31:0]);
			assign lsu_result_corr_r[31:0] = (((({32 {lsu_pkt_r[5] & lsu_pkt_r[11]}} & {24'b000000000000000000000000, lsu_ld_datafn_corr_r[7:0]}) | ({32 {lsu_pkt_r[5] & lsu_pkt_r[10]}} & {16'b0000000000000000, lsu_ld_datafn_corr_r[15:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[11]}} & {{24 {lsu_ld_datafn_corr_r[7]}}, lsu_ld_datafn_corr_r[7:0]})) | ({32 {~lsu_pkt_r[5] & lsu_pkt_r[10]}} & {{16 {lsu_ld_datafn_corr_r[15]}}, lsu_ld_datafn_corr_r[15:0]})) | ({32 {lsu_pkt_r[9]}} & lsu_ld_datafn_corr_r[31:0]);
		end
	endgenerate
	assign lsu_fir_addr[31:1] = lsu_ld_data_corr_r[31:1];
	assign lsu_addr_d[31:0] = full_addr_d[31:0];
	assign lsu_commit_r = ((lsu_pkt_r[0] & (lsu_pkt_r[6] | lsu_pkt_r[7])) & ~flush_r) & ~lsu_pkt_r[4];
	assign dma_mem_wdata_shifted[63:0] = dma_mem_wdata[63:0] >> {dma_mem_addr[2:0], 3'b000};
	assign store_data_d[31:0] = (dma_dccm_req ? dma_mem_wdata_shifted[31:0] : exu_lsu_rs2_d[31:0]);
	assign store_data_m_in[31:0] = (lsu_pkt_d[3] ? lsu_result_m[31:0] : store_data_d[31:0]);
	assign store_data_m[31:0] = (picm_mask_data_m[31:0] | {32 {~addr_in_pic_m}}) & (lsu_pkt_m[1] ? lsu_result_m[31:0] : store_data_pre_m[31:0]);
	rvdff #(.WIDTH(32)) sdmff(
		.rst_l(rst_l),
		.din(store_data_m_in[31:0]),
		.dout(store_data_pre_m[31:0]),
		.clk(lsu_store_c1_m_clk)
	);
	rvdff #(.WIDTH(32)) samff(
		.rst_l(rst_l),
		.din(lsu_addr_d[31:0]),
		.dout(lsu_addr_m[31:0]),
		.clk(lsu_c1_m_clk)
	);
	rvdff #(.WIDTH(32)) sarff(
		.rst_l(rst_l),
		.din(lsu_addr_m[31:0]),
		.dout(lsu_addr_r[31:0]),
		.clk(lsu_c1_r_clk)
	);
	assign end_addr_m[31:3] = (ldst_dual_m ? end_addr_pre_m[31:3] : lsu_addr_m[31:3]);
	assign end_addr_r[31:3] = (ldst_dual_r ? end_addr_pre_r[31:3] : lsu_addr_r[31:3]);
	rvdffe #(.WIDTH(29)) end_addr_hi_mff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(end_addr_d[31:3]),
		.dout(end_addr_pre_m[31:3]),
		.en((lsu_pkt_d[0] & ldst_dual_d) | clk_override)
	);
	rvdffe #(.WIDTH(29)) end_addr_hi_rff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(end_addr_m[31:3]),
		.dout(end_addr_pre_r[31:3]),
		.en((lsu_pkt_m[0] & ldst_dual_m) | clk_override)
	);
	rvdff #(.WIDTH(3)) end_addr_lo_mff(
		.rst_l(rst_l),
		.din(end_addr_d[2:0]),
		.dout(end_addr_m[2:0]),
		.clk(lsu_c1_m_clk)
	);
	rvdff #(.WIDTH(3)) end_addr_lo_rff(
		.rst_l(rst_l),
		.din(end_addr_m[2:0]),
		.dout(end_addr_r[2:0]),
		.clk(lsu_c1_r_clk)
	);
	rvdff #(.WIDTH(1)) addr_in_dccm_mff(
		.din(addr_in_dccm_d),
		.dout(addr_in_dccm_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) addr_in_dccm_rff(
		.din(addr_in_dccm_m),
		.dout(addr_in_dccm_r),
		.clk(lsu_c1_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) addr_in_pic_mff(
		.din(addr_in_pic_d),
		.dout(addr_in_pic_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) addr_in_pic_rff(
		.din(addr_in_pic_m),
		.dout(addr_in_pic_r),
		.clk(lsu_c1_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) addr_external_mff(
		.din(addr_external_d),
		.dout(addr_external_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) addr_external_rff(
		.din(addr_external_m),
		.dout(addr_external_r),
		.clk(lsu_c1_r_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) access_fault_mff(
		.din(access_fault_d),
		.dout(access_fault_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) misaligned_fault_mff(
		.din(misaligned_fault_d),
		.dout(misaligned_fault_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(4)) exc_mscause_mff(
		.din(exc_mscause_d[3:0]),
		.dout(exc_mscause_m[3:0]),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) fir_dccm_access_error_mff(
		.din(fir_dccm_access_error_d),
		.dout(fir_dccm_access_error_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdff #(.WIDTH(1)) fir_nondccm_access_error_mff(
		.din(fir_nondccm_access_error_d),
		.dout(fir_nondccm_access_error_m),
		.clk(lsu_c1_m_clk),
		.rst_l(rst_l)
	);
	rvdffe #(.WIDTH(32)) bus_read_data_r_ff(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(bus_read_data_m[31:0]),
		.dout(bus_read_data_r[31:0]),
		.en(addr_external_m | clk_override)
	);
endmodule
module eb1_lsu_stbuf (
	clk,
	rst_l,
	lsu_stbuf_c1_clk,
	lsu_free_c2_clk,
	store_stbuf_reqvld_r,
	lsu_commit_r,
	dec_lsu_valid_raw_d,
	store_data_hi_r,
	store_data_lo_r,
	store_datafn_hi_r,
	store_datafn_lo_r,
	stbuf_reqvld_any,
	stbuf_reqvld_flushed_any,
	stbuf_addr_any,
	stbuf_data_any,
	lsu_stbuf_commit_any,
	lsu_stbuf_full_any,
	lsu_stbuf_empty_any,
	ldst_stbuf_reqvld_r,
	lsu_addr_d,
	lsu_addr_m,
	lsu_addr_r,
	end_addr_d,
	end_addr_m,
	end_addr_r,
	ldst_dual_d,
	ldst_dual_m,
	ldst_dual_r,
	addr_in_dccm_m,
	addr_in_dccm_r,
	lsu_cmpen_m,
	lsu_pkt_m,
	lsu_pkt_r,
	stbuf_fwddata_hi_m,
	stbuf_fwddata_lo_m,
	stbuf_fwdbyteen_hi_m,
	stbuf_fwdbyteen_lo_m,
	scan_mode
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire clk;
	input wire rst_l;
	input wire lsu_stbuf_c1_clk;
	input wire lsu_free_c2_clk;
	input wire store_stbuf_reqvld_r;
	input wire lsu_commit_r;
	input wire dec_lsu_valid_raw_d;
	input wire [pt[1382-:10] - 1:0] store_data_hi_r;
	input wire [pt[1382-:10] - 1:0] store_data_lo_r;
	input wire [pt[1382-:10] - 1:0] store_datafn_hi_r;
	input wire [pt[1382-:10] - 1:0] store_datafn_lo_r;
	output wire stbuf_reqvld_any;
	output wire stbuf_reqvld_flushed_any;
	output wire [pt[157-:9] - 1:0] stbuf_addr_any;
	output wire [pt[1382-:10] - 1:0] stbuf_data_any;
	input wire lsu_stbuf_commit_any;
	output wire lsu_stbuf_full_any;
	output wire lsu_stbuf_empty_any;
	output wire ldst_stbuf_reqvld_r;
	input wire [pt[157-:9] - 1:0] lsu_addr_d;
	input wire [31:0] lsu_addr_m;
	input wire [31:0] lsu_addr_r;
	input wire [pt[157-:9] - 1:0] end_addr_d;
	input wire [31:0] end_addr_m;
	input wire [31:0] end_addr_r;
	input wire ldst_dual_d;
	input wire ldst_dual_m;
	input wire ldst_dual_r;
	input wire addr_in_dccm_m;
	input wire addr_in_dccm_r;
	input wire lsu_cmpen_m;
	input wire [13:0] lsu_pkt_m;
	input wire [13:0] lsu_pkt_r;
	output wire [pt[1382-:10] - 1:0] stbuf_fwddata_hi_m;
	output wire [pt[1382-:10] - 1:0] stbuf_fwddata_lo_m;
	output wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_hi_m;
	output wire [pt[1389-:7] - 1:0] stbuf_fwdbyteen_lo_m;
	input wire scan_mode;
	localparam DEPTH = pt[148-:8];
	localparam DATA_WIDTH = pt[1382-:10];
	localparam BYTE_WIDTH = pt[1389-:7];
	localparam DEPTH_LOG2 = $clog2(DEPTH);
	wire [DEPTH - 1:0] stbuf_vld;
	wire [DEPTH - 1:0] stbuf_dma_kill;
	wire [(DEPTH * pt[157-:9]) - 1:0] stbuf_addr;
	wire [(DEPTH * BYTE_WIDTH) - 1:0] stbuf_byteen;
	wire [(DEPTH * DATA_WIDTH) - 1:0] stbuf_data;
	wire [DEPTH - 1:0] sel_lo;
	wire [DEPTH - 1:0] stbuf_wr_en;
	reg [DEPTH - 1:0] stbuf_dma_kill_en;
	wire [DEPTH - 1:0] stbuf_reset;
	wire [(DEPTH * pt[157-:9]) - 1:0] stbuf_addrin;
	wire [(DEPTH * DATA_WIDTH) - 1:0] stbuf_datain;
	wire [(DEPTH * BYTE_WIDTH) - 1:0] stbuf_byteenin;
	wire [7:0] store_byteen_ext_r;
	wire [BYTE_WIDTH - 1:0] store_byteen_hi_r;
	wire [BYTE_WIDTH - 1:0] store_byteen_lo_r;
	wire WrPtrEn;
	wire RdPtrEn;
	wire [DEPTH_LOG2 - 1:0] WrPtr;
	wire [DEPTH_LOG2 - 1:0] RdPtr;
	wire [DEPTH_LOG2 - 1:0] NxtWrPtr;
	wire [DEPTH_LOG2 - 1:0] NxtRdPtr;
	wire [DEPTH_LOG2 - 1:0] WrPtrPlus1;
	wire [DEPTH_LOG2 - 1:0] WrPtrPlus2;
	wire [DEPTH_LOG2 - 1:0] RdPtrPlus1;
	wire dual_stbuf_write_r;
	wire isdccmst_m;
	wire isdccmst_r;
	reg [3:0] stbuf_numvld_any;
	wire [3:0] stbuf_specvld_any;
	wire [1:0] stbuf_specvld_m;
	wire [1:0] stbuf_specvld_r;
	wire [pt[157-:9] - 1:$clog2(BYTE_WIDTH)] cmpaddr_hi_m;
	wire [pt[157-:9] - 1:$clog2(BYTE_WIDTH)] cmpaddr_lo_m;
	reg [DEPTH - 1:0] stbuf_match_hi;
	reg [DEPTH - 1:0] stbuf_match_lo;
	reg [(DEPTH * BYTE_WIDTH) - 1:0] stbuf_fwdbyteenvec_hi;
	reg [(DEPTH * BYTE_WIDTH) - 1:0] stbuf_fwdbyteenvec_lo;
	reg [DATA_WIDTH - 1:0] stbuf_fwddata_hi_pre_m;
	reg [DATA_WIDTH - 1:0] stbuf_fwddata_lo_pre_m;
	reg [BYTE_WIDTH - 1:0] stbuf_fwdbyteen_hi_pre_m;
	reg [BYTE_WIDTH - 1:0] stbuf_fwdbyteen_lo_pre_m;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_lo_lo;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_hi_lo;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_lo_hi;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_hi_hi;
	wire ld_addr_rhit_lo_lo;
	wire ld_addr_rhit_hi_lo;
	wire ld_addr_rhit_lo_hi;
	wire ld_addr_rhit_hi_hi;
	wire [BYTE_WIDTH - 1:0] ld_byte_hit_lo;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_lo;
	wire [BYTE_WIDTH - 1:0] ld_byte_hit_hi;
	wire [BYTE_WIDTH - 1:0] ld_byte_rhit_hi;
	wire [BYTE_WIDTH - 1:0] ldst_byteen_hi_r;
	wire [BYTE_WIDTH - 1:0] ldst_byteen_lo_r;
	wire [7:0] ldst_byteen_r;
	wire [7:0] ldst_byteen_ext_r;
	wire [31:0] ld_fwddata_rpipe_lo;
	wire [31:0] ld_fwddata_rpipe_hi;
	wire [DEPTH - 1:0] store_matchvec_lo_r;
	wire [DEPTH - 1:0] store_matchvec_hi_r;
	wire store_coalesce_lo_r;
	wire store_coalesce_hi_r;
	assign store_byteen_ext_r[7:0] = ldst_byteen_r[7:0] << lsu_addr_r[1:0];
	assign store_byteen_hi_r[BYTE_WIDTH - 1:0] = store_byteen_ext_r[7:4] & {4 {lsu_pkt_r[6]}};
	assign store_byteen_lo_r[BYTE_WIDTH - 1:0] = store_byteen_ext_r[3:0] & {4 {lsu_pkt_r[6]}};
	assign RdPtrPlus1[DEPTH_LOG2 - 1:0] = RdPtr[DEPTH_LOG2 - 1:0] + 1'b1;
	assign WrPtrPlus1[DEPTH_LOG2 - 1:0] = WrPtr[DEPTH_LOG2 - 1:0] + 1'b1;
	assign WrPtrPlus2[DEPTH_LOG2 - 1:0] = WrPtr[DEPTH_LOG2 - 1:0] + 2'b10;
	assign dual_stbuf_write_r = ldst_dual_r & store_stbuf_reqvld_r;
	assign ldst_stbuf_reqvld_r = (lsu_commit_r | lsu_pkt_r[4]) & store_stbuf_reqvld_r;
	generate
		genvar i;
		for (i = 0; i < DEPTH; i = i + 1) begin : FindMatchEntry
			assign store_matchvec_lo_r[i] = (((stbuf_addr[(i * pt[157-:9]) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? pt[157-:9] - 1 : ((pt[157-:9] - 1) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)) - 1)-:((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)] == lsu_addr_r[pt[157-:9] - 1:$clog2(BYTE_WIDTH)]) & stbuf_vld[i]) & ~stbuf_dma_kill[i]) & ~stbuf_reset[i];
			assign store_matchvec_hi_r[i] = ((((stbuf_addr[(i * pt[157-:9]) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? pt[157-:9] - 1 : ((pt[157-:9] - 1) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)) - 1)-:((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)] == end_addr_r[pt[157-:9] - 1:$clog2(BYTE_WIDTH)]) & stbuf_vld[i]) & ~stbuf_dma_kill[i]) & dual_stbuf_write_r) & ~stbuf_reset[i];
		end
	endgenerate
	assign store_coalesce_lo_r = |store_matchvec_lo_r[DEPTH - 1:0];
	assign store_coalesce_hi_r = |store_matchvec_hi_r[DEPTH - 1:0];
	generate
		if (pt[1365-:5] == 1) begin : Gen_dccm_enable
			for (i = 0; i < DEPTH; i = i + 1) begin : GenStBuf
				assign stbuf_wr_en[i] = ldst_stbuf_reqvld_r & ((((((i == WrPtr[DEPTH_LOG2 - 1:0]) & ~store_coalesce_lo_r) | (((i == WrPtr[DEPTH_LOG2 - 1:0]) & dual_stbuf_write_r) & ~store_coalesce_hi_r)) | (((i == WrPtrPlus1[DEPTH_LOG2 - 1:0]) & dual_stbuf_write_r) & ~(store_coalesce_lo_r | store_coalesce_hi_r))) | store_matchvec_lo_r[i]) | store_matchvec_hi_r[i]);
				assign stbuf_reset[i] = (lsu_stbuf_commit_any | stbuf_reqvld_flushed_any) & (i == RdPtr[DEPTH_LOG2 - 1:0]);
				assign sel_lo[i] = (((~ldst_dual_r | store_stbuf_reqvld_r) & (i == WrPtr[DEPTH_LOG2 - 1:0])) & ~store_coalesce_lo_r) | store_matchvec_lo_r[i];
				assign stbuf_addrin[(i * pt[157-:9]) + (pt[157-:9] - 1)-:pt[157-:9]] = (sel_lo[i] ? lsu_addr_r[pt[157-:9] - 1:0] : end_addr_r[pt[157-:9] - 1:0]);
				assign stbuf_byteenin[(i * BYTE_WIDTH) + (BYTE_WIDTH - 1)-:BYTE_WIDTH] = (sel_lo[i] ? stbuf_byteen[(i * BYTE_WIDTH) + (BYTE_WIDTH - 1)-:BYTE_WIDTH] | store_byteen_lo_r[BYTE_WIDTH - 1:0] : stbuf_byteen[(i * BYTE_WIDTH) + (BYTE_WIDTH - 1)-:BYTE_WIDTH] | store_byteen_hi_r[BYTE_WIDTH - 1:0]);
				assign stbuf_datain[(i * DATA_WIDTH) + 7-:8] = (sel_lo[i] ? (~stbuf_byteen[i * BYTE_WIDTH] | store_byteen_lo_r[0] ? store_datafn_lo_r[7:0] : stbuf_data[(i * DATA_WIDTH) + 7-:8]) : (~stbuf_byteen[i * BYTE_WIDTH] | store_byteen_hi_r[0] ? store_datafn_hi_r[7:0] : stbuf_data[(i * DATA_WIDTH) + 7-:8]));
				assign stbuf_datain[(i * DATA_WIDTH) + 15-:8] = (sel_lo[i] ? (~stbuf_byteen[(i * BYTE_WIDTH) + 1] | store_byteen_lo_r[1] ? store_datafn_lo_r[15:8] : stbuf_data[(i * DATA_WIDTH) + 15-:8]) : (~stbuf_byteen[(i * BYTE_WIDTH) + 1] | store_byteen_hi_r[1] ? store_datafn_hi_r[15:8] : stbuf_data[(i * DATA_WIDTH) + 15-:8]));
				assign stbuf_datain[(i * DATA_WIDTH) + 23-:8] = (sel_lo[i] ? (~stbuf_byteen[(i * BYTE_WIDTH) + 2] | store_byteen_lo_r[2] ? store_datafn_lo_r[23:16] : stbuf_data[(i * DATA_WIDTH) + 23-:8]) : (~stbuf_byteen[(i * BYTE_WIDTH) + 2] | store_byteen_hi_r[2] ? store_datafn_hi_r[23:16] : stbuf_data[(i * DATA_WIDTH) + 23-:8]));
				assign stbuf_datain[(i * DATA_WIDTH) + 31-:8] = (sel_lo[i] ? (~stbuf_byteen[(i * BYTE_WIDTH) + 3] | store_byteen_lo_r[3] ? store_datafn_lo_r[31:24] : stbuf_data[(i * DATA_WIDTH) + 31-:8]) : (~stbuf_byteen[(i * BYTE_WIDTH) + 3] | store_byteen_hi_r[3] ? store_datafn_hi_r[31:24] : stbuf_data[(i * DATA_WIDTH) + 31-:8]));
				rvdffsc #(.WIDTH(1)) stbuf_vldff(
					.din(1'b1),
					.dout(stbuf_vld[i]),
					.en(stbuf_wr_en[i]),
					.clear(stbuf_reset[i]),
					.clk(lsu_free_c2_clk),
					.rst_l(rst_l)
				);
				rvdffsc #(.WIDTH(1)) stbuf_killff(
					.din(1'b1),
					.dout(stbuf_dma_kill[i]),
					.en(stbuf_dma_kill_en[i]),
					.clear(stbuf_reset[i]),
					.clk(lsu_free_c2_clk),
					.rst_l(rst_l)
				);
				rvdffe #(.WIDTH(pt[157-:9])) stbuf_addrff(
					.din(stbuf_addrin[(i * pt[157-:9]) + (pt[157-:9] - 1)-:pt[157-:9]]),
					.dout(stbuf_addr[(i * pt[157-:9]) + (pt[157-:9] - 1)-:pt[157-:9]]),
					.en(stbuf_wr_en[i]),
					.clk(clk),
					.rst_l(rst_l),
					.scan_mode(scan_mode)
				);
				rvdffsc #(.WIDTH(BYTE_WIDTH)) stbuf_byteenff(
					.din(stbuf_byteenin[(i * BYTE_WIDTH) + (BYTE_WIDTH - 1)-:BYTE_WIDTH]),
					.dout(stbuf_byteen[(i * BYTE_WIDTH) + (BYTE_WIDTH - 1)-:BYTE_WIDTH]),
					.en(stbuf_wr_en[i]),
					.clear(stbuf_reset[i]),
					.clk(lsu_stbuf_c1_clk),
					.rst_l(rst_l)
				);
				rvdffe #(.WIDTH(DATA_WIDTH)) stbuf_dataff(
					.din(stbuf_datain[(i * DATA_WIDTH) + (DATA_WIDTH - 1)-:DATA_WIDTH]),
					.dout(stbuf_data[(i * DATA_WIDTH) + (DATA_WIDTH - 1)-:DATA_WIDTH]),
					.en(stbuf_wr_en[i]),
					.clk(clk),
					.rst_l(rst_l),
					.scan_mode(scan_mode)
				);
			end
		end
		else begin : Gen_dccm_disable
			assign stbuf_wr_en[DEPTH - 1:0] = {DEPTH {1'sb0}};
			assign stbuf_reset[DEPTH - 1:0] = {DEPTH {1'sb0}};
			assign stbuf_vld[DEPTH - 1:0] = {DEPTH {1'sb0}};
			assign stbuf_dma_kill[DEPTH - 1:0] = {DEPTH {1'sb0}};
			assign stbuf_addr[pt[157-:9] * ((DEPTH - 1) - (DEPTH - 1))+:pt[157-:9] * DEPTH] = {pt[157-:9] * DEPTH {1'sb0}};
			assign stbuf_byteen[BYTE_WIDTH * ((DEPTH - 1) - (DEPTH - 1))+:BYTE_WIDTH * DEPTH] = {BYTE_WIDTH * DEPTH {1'sb0}};
			assign stbuf_data[DATA_WIDTH * ((DEPTH - 1) - (DEPTH - 1))+:DATA_WIDTH * DEPTH] = {DATA_WIDTH * DEPTH {1'sb0}};
		end
	endgenerate
	assign stbuf_reqvld_flushed_any = stbuf_vld[RdPtr] & stbuf_dma_kill[RdPtr];
	assign stbuf_reqvld_any = (stbuf_vld[RdPtr] & ~stbuf_dma_kill[RdPtr]) & ~(|stbuf_dma_kill_en[DEPTH - 1:0]);
	assign stbuf_addr_any[pt[157-:9] - 1:0] = stbuf_addr[(RdPtr * pt[157-:9]) + (pt[157-:9] - 1)-:pt[157-:9]];
	assign stbuf_data_any[DATA_WIDTH - 1:0] = stbuf_data[(RdPtr * DATA_WIDTH) + (DATA_WIDTH - 1)-:DATA_WIDTH];
	assign WrPtrEn = ((ldst_stbuf_reqvld_r & ~dual_stbuf_write_r) & ~(store_coalesce_hi_r | store_coalesce_lo_r)) | ((ldst_stbuf_reqvld_r & dual_stbuf_write_r) & ~(store_coalesce_hi_r & store_coalesce_lo_r));
	assign NxtWrPtr[DEPTH_LOG2 - 1:0] = ((ldst_stbuf_reqvld_r & dual_stbuf_write_r) & ~(store_coalesce_hi_r | store_coalesce_lo_r) ? WrPtrPlus2[DEPTH_LOG2 - 1:0] : WrPtrPlus1[DEPTH_LOG2 - 1:0]);
	assign RdPtrEn = lsu_stbuf_commit_any | stbuf_reqvld_flushed_any;
	assign NxtRdPtr[DEPTH_LOG2 - 1:0] = RdPtrPlus1[DEPTH_LOG2 - 1:0];
	always @(*) begin
		stbuf_numvld_any[3:0] = {4 {1'sb0}};
		begin : sv2v_autoblock_59
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				stbuf_numvld_any[3:0] = stbuf_numvld_any[3:0] + {3'b000, stbuf_vld[i]};
		end
	end
	assign isdccmst_m = ((lsu_pkt_m[0] & lsu_pkt_m[6]) & addr_in_dccm_m) & ~lsu_pkt_m[4];
	assign isdccmst_r = ((lsu_pkt_r[0] & lsu_pkt_r[6]) & addr_in_dccm_r) & ~lsu_pkt_r[4];
	assign stbuf_specvld_m[1:0] = {1'b0, isdccmst_m} << (isdccmst_m & ldst_dual_m);
	assign stbuf_specvld_r[1:0] = {1'b0, isdccmst_r} << (isdccmst_r & ldst_dual_r);
	assign stbuf_specvld_any[3:0] = (stbuf_numvld_any[3:0] + {2'b00, stbuf_specvld_m[1:0]}) + {2'b00, stbuf_specvld_r[1:0]};
	assign lsu_stbuf_full_any = (~ldst_dual_d & dec_lsu_valid_raw_d ? stbuf_specvld_any[3:0] >= DEPTH : stbuf_specvld_any[3:0] >= (DEPTH - 1));
	assign lsu_stbuf_empty_any = stbuf_numvld_any[3:0] == 4'b0000;
	assign cmpaddr_hi_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)] = end_addr_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)];
	assign cmpaddr_lo_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)] = lsu_addr_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)];
	always @(*) begin : GenLdFwd
		stbuf_fwdbyteen_hi_pre_m[BYTE_WIDTH - 1:0] = {BYTE_WIDTH {1'sb0}};
		stbuf_fwdbyteen_lo_pre_m[BYTE_WIDTH - 1:0] = {BYTE_WIDTH {1'sb0}};
		begin : sv2v_autoblock_60
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					stbuf_match_hi[i] = (((stbuf_addr[(i * pt[157-:9]) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? pt[157-:9] - 1 : ((pt[157-:9] - 1) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)) - 1)-:((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)] == cmpaddr_hi_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)]) & stbuf_vld[i]) & ~stbuf_dma_kill[i]) & addr_in_dccm_m;
					stbuf_match_lo[i] = (((stbuf_addr[(i * pt[157-:9]) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? pt[157-:9] - 1 : ((pt[157-:9] - 1) + ((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)) - 1)-:((pt[157-:9] - 1) >= $clog2(BYTE_WIDTH) ? ((pt[157-:9] - 1) - $clog2(BYTE_WIDTH)) + 1 : ($clog2(BYTE_WIDTH) - (pt[157-:9] - 1)) + 1)] == cmpaddr_lo_m[pt[157-:9] - 1:$clog2(BYTE_WIDTH)]) & stbuf_vld[i]) & ~stbuf_dma_kill[i]) & addr_in_dccm_m;
					stbuf_dma_kill_en[i] = (((stbuf_match_hi[i] | stbuf_match_lo[i]) & lsu_pkt_m[0]) & lsu_pkt_m[4]) & lsu_pkt_m[6];
					begin : sv2v_autoblock_61
						reg signed [31:0] j;
						for (j = 0; j < BYTE_WIDTH; j = j + 1)
							begin
								stbuf_fwdbyteenvec_hi[(i * BYTE_WIDTH) + j] = (stbuf_match_hi[i] & stbuf_byteen[(i * BYTE_WIDTH) + j]) & stbuf_vld[i];
								stbuf_fwdbyteen_hi_pre_m[j] = stbuf_fwdbyteen_hi_pre_m[j] | stbuf_fwdbyteenvec_hi[(i * BYTE_WIDTH) + j];
								stbuf_fwdbyteenvec_lo[(i * BYTE_WIDTH) + j] = (stbuf_match_lo[i] & stbuf_byteen[(i * BYTE_WIDTH) + j]) & stbuf_vld[i];
								stbuf_fwdbyteen_lo_pre_m[j] = stbuf_fwdbyteen_lo_pre_m[j] | stbuf_fwdbyteenvec_lo[(i * BYTE_WIDTH) + j];
							end
					end
				end
		end
	end
	always @(*) begin : GenLdData
		stbuf_fwddata_hi_pre_m[31:0] = {32 {1'sb0}};
		stbuf_fwddata_lo_pre_m[31:0] = {32 {1'sb0}};
		begin : sv2v_autoblock_62
			reg signed [31:0] i;
			for (i = 0; i < DEPTH; i = i + 1)
				begin
					stbuf_fwddata_hi_pre_m[31:0] = stbuf_fwddata_hi_pre_m[31:0] | ({32 {stbuf_match_hi[i]}} & stbuf_data[(i * DATA_WIDTH) + 31-:32]);
					stbuf_fwddata_lo_pre_m[31:0] = stbuf_fwddata_lo_pre_m[31:0] | ({32 {stbuf_match_lo[i]}} & stbuf_data[(i * DATA_WIDTH) + 31-:32]);
				end
		end
	end
	assign ldst_byteen_r[7:0] = ((({8 {lsu_pkt_r[11]}} & 8'b00000001) | ({8 {lsu_pkt_r[10]}} & 8'b00000011)) | ({8 {lsu_pkt_r[9]}} & 8'b00001111)) | ({8 {lsu_pkt_r[8]}} & 8'b11111111);
	assign ldst_byteen_ext_r[7:0] = ldst_byteen_r[7:0] << lsu_addr_r[1:0];
	assign ldst_byteen_hi_r[3:0] = ldst_byteen_ext_r[7:4];
	assign ldst_byteen_lo_r[3:0] = ldst_byteen_ext_r[3:0];
	assign ld_addr_rhit_lo_lo = (((lsu_addr_m[31:2] == lsu_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & ~lsu_pkt_r[4];
	assign ld_addr_rhit_lo_hi = (((end_addr_m[31:2] == lsu_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & ~lsu_pkt_r[4];
	assign ld_addr_rhit_hi_lo = ((((lsu_addr_m[31:2] == end_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & ~lsu_pkt_r[4]) & dual_stbuf_write_r;
	assign ld_addr_rhit_hi_hi = ((((end_addr_m[31:2] == end_addr_r[31:2]) & lsu_pkt_r[0]) & lsu_pkt_r[6]) & ~lsu_pkt_r[4]) & dual_stbuf_write_r;
	generate
		for (i = 0; i < BYTE_WIDTH; i = i + 1) begin
			assign ld_byte_rhit_lo_lo[i] = ld_addr_rhit_lo_lo & ldst_byteen_lo_r[i];
			assign ld_byte_rhit_lo_hi[i] = ld_addr_rhit_lo_hi & ldst_byteen_lo_r[i];
			assign ld_byte_rhit_hi_lo[i] = ld_addr_rhit_hi_lo & ldst_byteen_hi_r[i];
			assign ld_byte_rhit_hi_hi[i] = ld_addr_rhit_hi_hi & ldst_byteen_hi_r[i];
			assign ld_byte_rhit_lo[i] = ld_byte_rhit_lo_lo[i] | ld_byte_rhit_hi_lo[i];
			assign ld_byte_rhit_hi[i] = ld_byte_rhit_lo_hi[i] | ld_byte_rhit_hi_hi[i];
			assign ld_fwddata_rpipe_lo[(8 * i) + 7:8 * i] = ({8 {ld_byte_rhit_lo_lo[i]}} & store_data_lo_r[(8 * i) + 7:8 * i]) | ({8 {ld_byte_rhit_hi_lo[i]}} & store_data_hi_r[(8 * i) + 7:8 * i]);
			assign ld_fwddata_rpipe_hi[(8 * i) + 7:8 * i] = ({8 {ld_byte_rhit_lo_hi[i]}} & store_data_lo_r[(8 * i) + 7:8 * i]) | ({8 {ld_byte_rhit_hi_hi[i]}} & store_data_hi_r[(8 * i) + 7:8 * i]);
			assign ld_byte_hit_lo[i] = ld_byte_rhit_lo_lo[i] | ld_byte_rhit_hi_lo[i];
			assign ld_byte_hit_hi[i] = ld_byte_rhit_lo_hi[i] | ld_byte_rhit_hi_hi[i];
			assign stbuf_fwdbyteen_hi_m[i] = ld_byte_hit_hi[i] | stbuf_fwdbyteen_hi_pre_m[i];
			assign stbuf_fwdbyteen_lo_m[i] = ld_byte_hit_lo[i] | stbuf_fwdbyteen_lo_pre_m[i];
			assign stbuf_fwddata_lo_m[(8 * i) + 7:8 * i] = (ld_byte_rhit_lo[i] ? ld_fwddata_rpipe_lo[(8 * i) + 7:8 * i] : stbuf_fwddata_lo_pre_m[(8 * i) + 7:8 * i]);
			assign stbuf_fwddata_hi_m[(8 * i) + 7:8 * i] = (ld_byte_rhit_hi[i] ? ld_fwddata_rpipe_hi[(8 * i) + 7:8 * i] : stbuf_fwddata_hi_pre_m[(8 * i) + 7:8 * i]);
		end
	endgenerate
	rvdffs #(.WIDTH(DEPTH_LOG2)) WrPtrff(
		.din(NxtWrPtr[DEPTH_LOG2 - 1:0]),
		.dout(WrPtr[DEPTH_LOG2 - 1:0]),
		.en(WrPtrEn),
		.clk(lsu_stbuf_c1_clk),
		.rst_l(rst_l)
	);
	rvdffs #(.WIDTH(DEPTH_LOG2)) RdPtrff(
		.din(NxtRdPtr[DEPTH_LOG2 - 1:0]),
		.dout(RdPtr[DEPTH_LOG2 - 1:0]),
		.en(RdPtrEn),
		.clk(lsu_stbuf_c1_clk),
		.rst_l(rst_l)
	);
endmodule
module eb1_lsu_trigger (
	trigger_pkt_any,
	lsu_pkt_m,
	lsu_addr_m,
	store_data_m,
	lsu_trigger_match_m
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [151:0] trigger_pkt_any;
	input wire [13:0] lsu_pkt_m;
	input wire [31:0] lsu_addr_m;
	input wire [31:0] store_data_m;
	output wire [3:0] lsu_trigger_match_m;
	reg trigger_enable;
	wire [127:0] lsu_match_data;
	wire [3:0] lsu_trigger_data_match;
	wire [31:0] store_data_trigger_m;
	wire [31:0] ldst_addr_trigger_m;
	always @(*) begin
		trigger_enable = 1'b0;
		begin : sv2v_autoblock_63
			reg signed [31:0] i;
			for (i = 0; i < 4; i = i + 1)
				trigger_enable = trigger_enable | trigger_pkt_any[(i * 38) + 32];
		end
	end
	assign store_data_trigger_m[31:0] = {{16 {lsu_pkt_m[9]}} & store_data_m[31:16], {8 {lsu_pkt_m[10] | lsu_pkt_m[9]}} & store_data_m[15:8], store_data_m[7:0]} & {32 {trigger_enable}};
	assign ldst_addr_trigger_m[31:0] = lsu_addr_m[31:0] & {32 {trigger_enable}};
	generate
		genvar i;
		for (i = 0; i < 4; i = i + 1) begin
			assign lsu_match_data[(i * 32) + 31-:32] = ({32 {~trigger_pkt_any[(i * 38) + 37]}} & ldst_addr_trigger_m[31:0]) | ({32 {trigger_pkt_any[(i * 38) + 37] & trigger_pkt_any[(i * 38) + 35]}} & store_data_trigger_m[31:0]);
			rvmaskandmatch trigger_match(
				.mask(trigger_pkt_any[(i * 38) + 31-:32]),
				.data(lsu_match_data[(i * 32) + 31-:32]),
				.masken(trigger_pkt_any[(i * 38) + 36]),
				.match(lsu_trigger_data_match[i])
			);
			assign lsu_trigger_match_m[i] = (((lsu_pkt_m[0] & ~lsu_pkt_m[4]) & trigger_enable) & ((trigger_pkt_any[(i * 38) + 35] & lsu_pkt_m[6]) | ((trigger_pkt_any[(i * 38) + 34] & lsu_pkt_m[7]) & ~trigger_pkt_any[(i * 38) + 37]))) & lsu_trigger_data_match[i];
		end
	endgenerate
endmodule
module rvjtag_tap (
	trst,
	tck,
	tms,
	tdi,
	tdo,
	tdoEnable,
	wr_data,
	wr_addr,
	wr_en,
	rd_en,
	rd_data,
	rd_status,
	dmi_reset,
	dmi_hard_reset,
	idle,
	dmi_stat,
	jtag_id,
	version
);
	parameter AWIDTH = 7;
	input trst;
	input tck;
	input tms;
	input tdi;
	output reg tdo;
	output tdoEnable;
	output [31:0] wr_data;
	output [AWIDTH - 1:0] wr_addr;
	output wr_en;
	output rd_en;
	input [31:0] rd_data;
	input [1:0] rd_status;
	output reg dmi_reset;
	output reg dmi_hard_reset;
	input [2:0] idle;
	input [1:0] dmi_stat;
	input [31:1] jtag_id;
	input [3:0] version;
	localparam USER_DR_LENGTH = AWIDTH + 34;
	reg [USER_DR_LENGTH - 1:0] sr;
	reg [USER_DR_LENGTH - 1:0] nsr;
	reg [USER_DR_LENGTH - 1:0] dr;
	reg [3:0] state;
	reg [3:0] nstate;
	reg [4:0] ir;
	wire jtag_reset;
	wire shift_dr;
	wire pause_dr;
	wire update_dr;
	wire capture_dr;
	wire shift_ir;
	wire pause_ir;
	wire update_ir;
	wire capture_ir;
	wire [1:0] dr_en;
	wire devid_sel;
	wire [5:0] abits;
	assign abits = AWIDTH[5:0];
	localparam TEST_LOGIC_RESET_STATE = 0;
	localparam RUN_TEST_IDLE_STATE = 1;
	localparam SELECT_DR_SCAN_STATE = 2;
	localparam CAPTURE_DR_STATE = 3;
	localparam SHIFT_DR_STATE = 4;
	localparam EXIT1_DR_STATE = 5;
	localparam PAUSE_DR_STATE = 6;
	localparam EXIT2_DR_STATE = 7;
	localparam UPDATE_DR_STATE = 8;
	localparam SELECT_IR_SCAN_STATE = 9;
	localparam CAPTURE_IR_STATE = 10;
	localparam SHIFT_IR_STATE = 11;
	localparam EXIT1_IR_STATE = 12;
	localparam PAUSE_IR_STATE = 13;
	localparam EXIT2_IR_STATE = 14;
	localparam UPDATE_IR_STATE = 15;
	always @(*) begin
		nstate = state;
		case (state)
			TEST_LOGIC_RESET_STATE: nstate = (tms ? TEST_LOGIC_RESET_STATE : RUN_TEST_IDLE_STATE);
			RUN_TEST_IDLE_STATE: nstate = (tms ? SELECT_DR_SCAN_STATE : RUN_TEST_IDLE_STATE);
			SELECT_DR_SCAN_STATE: nstate = (tms ? SELECT_IR_SCAN_STATE : CAPTURE_DR_STATE);
			CAPTURE_DR_STATE: nstate = (tms ? EXIT1_DR_STATE : SHIFT_DR_STATE);
			SHIFT_DR_STATE: nstate = (tms ? EXIT1_DR_STATE : SHIFT_DR_STATE);
			EXIT1_DR_STATE: nstate = (tms ? UPDATE_DR_STATE : PAUSE_DR_STATE);
			PAUSE_DR_STATE: nstate = (tms ? EXIT2_DR_STATE : PAUSE_DR_STATE);
			EXIT2_DR_STATE: nstate = (tms ? UPDATE_DR_STATE : SHIFT_DR_STATE);
			UPDATE_DR_STATE: nstate = (tms ? SELECT_DR_SCAN_STATE : RUN_TEST_IDLE_STATE);
			SELECT_IR_SCAN_STATE: nstate = (tms ? TEST_LOGIC_RESET_STATE : CAPTURE_IR_STATE);
			CAPTURE_IR_STATE: nstate = (tms ? EXIT1_IR_STATE : SHIFT_IR_STATE);
			SHIFT_IR_STATE: nstate = (tms ? EXIT1_IR_STATE : SHIFT_IR_STATE);
			EXIT1_IR_STATE: nstate = (tms ? UPDATE_IR_STATE : PAUSE_IR_STATE);
			PAUSE_IR_STATE: nstate = (tms ? EXIT2_IR_STATE : PAUSE_IR_STATE);
			EXIT2_IR_STATE: nstate = (tms ? UPDATE_IR_STATE : SHIFT_IR_STATE);
			UPDATE_IR_STATE: nstate = (tms ? SELECT_DR_SCAN_STATE : RUN_TEST_IDLE_STATE);
			default: nstate = TEST_LOGIC_RESET_STATE;
		endcase
	end
	always @(posedge tck or negedge trst)
		if (!trst)
			state <= TEST_LOGIC_RESET_STATE;
		else
			state <= nstate;
	assign jtag_reset = state == TEST_LOGIC_RESET_STATE;
	assign shift_dr = state == SHIFT_DR_STATE;
	assign pause_dr = state == PAUSE_DR_STATE;
	assign update_dr = state == UPDATE_DR_STATE;
	assign capture_dr = state == CAPTURE_DR_STATE;
	assign shift_ir = state == SHIFT_IR_STATE;
	assign pause_ir = state == PAUSE_IR_STATE;
	assign update_ir = state == UPDATE_IR_STATE;
	assign capture_ir = state == CAPTURE_IR_STATE;
	assign tdoEnable = shift_dr | shift_ir;
	always @(negedge tck or negedge trst)
		if (!trst)
			ir <= 5'b00001;
		else if (jtag_reset)
			ir <= 5'b00001;
		else if (update_ir)
			ir <= (sr[4:0] == {5 {1'sb0}} ? 5'h1f : sr[4:0]);
	assign devid_sel = ir == 5'b00001;
	assign dr_en[0] = ir == 5'b10000;
	assign dr_en[1] = ir == 5'b10001;
	always @(posedge tck or negedge trst)
		if (!trst)
			sr <= {USER_DR_LENGTH {1'sb0}};
		else
			sr <= nsr;
	always @(*) begin
		nsr = sr;
		case (1)
			shift_dr:
				case (1)
					dr_en[1]: nsr = {tdi, sr[USER_DR_LENGTH - 1:1]};
					dr_en[0], devid_sel: nsr = {{USER_DR_LENGTH - 32 {1'b0}}, tdi, sr[31:1]};
					default: nsr = {{USER_DR_LENGTH - 1 {1'b0}}, tdi};
				endcase
			capture_dr: begin
				nsr[0] = 1'b0;
				case (1)
					dr_en[0]: nsr = {{USER_DR_LENGTH - 15 {1'b0}}, idle, dmi_stat, abits, version};
					dr_en[1]: nsr = {{AWIDTH {1'b0}}, rd_data, rd_status};
					devid_sel: nsr = {{USER_DR_LENGTH - 32 {1'b0}}, jtag_id, 1'b1};
				endcase
			end
			shift_ir: nsr = {{USER_DR_LENGTH - 5 {1'b0}}, tdi, sr[4:1]};
			capture_ir: nsr = {{USER_DR_LENGTH - 1 {1'b0}}, 1'b1};
		endcase
	end
	always @(negedge tck) tdo <= sr[0];
	always @(posedge tck or negedge trst)
		if (!trst) begin
			dmi_hard_reset <= 1'b0;
			dmi_reset <= 1'b0;
		end
		else if (update_dr & dr_en[0]) begin
			dmi_hard_reset <= sr[17];
			dmi_reset <= sr[16];
		end
		else begin
			dmi_hard_reset <= 1'b0;
			dmi_reset <= 1'b0;
		end
	always @(posedge tck or negedge trst)
		if (!trst)
			dr <= {USER_DR_LENGTH {1'sb0}};
		else if (update_dr & dr_en[1])
			dr <= sr;
		else
			dr <= {dr[USER_DR_LENGTH - 1:2], 2'b00};
	assign {wr_addr, wr_data, wr_en, rd_en} = dr;
endmodule
module eb1_btb_tag_hash (
	pc,
	hash
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1] pc;
	output wire [pt[2139-:9] - 1:0] hash;
	assign hash = {(pc[((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + pt[2139-:9]:((pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]) + 1] ^ pc[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:(pt[2172-:9] + pt[2139-:9]) + 1]) ^ pc[pt[2172-:9] + pt[2139-:9]:pt[2172-:9] + 1]};
endmodule
module eb1_btb_tag_hash_fold (
	pc,
	hash
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:pt[2172-:9] + 1] pc;
	output wire [pt[2139-:9] - 1:0] hash;
	assign hash = {pc[(pt[2172-:9] + pt[2139-:9]) + pt[2139-:9]:(pt[2172-:9] + pt[2139-:9]) + 1] ^ pc[pt[2172-:9] + pt[2139-:9]:pt[2172-:9] + 1]};
endmodule
module eb1_btb_addr_hash (
	pc,
	hash
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [pt[2079-:9]:pt[2106-:9]] pc;
	output wire [pt[2172-:9]:pt[2163-:6]] hash;
	generate
		if (pt[2125-:5]) begin : fold2
			assign hash[pt[2172-:9]:pt[2163-:6]] = pc[pt[2115-:9]:pt[2106-:9]] ^ pc[pt[2079-:9]:pt[2070-:9]];
		end
		else assign hash[pt[2172-:9]:pt[2163-:6]] = (pc[pt[2115-:9]:pt[2106-:9]] ^ pc[pt[2097-:9]:pt[2088-:9]]) ^ pc[pt[2079-:9]:pt[2070-:9]];
	endgenerate
endmodule
module eb1_btb_ghr_hash (
	hashin,
	ghr,
	hash
);
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	parameter [2270:0] pt = {232'h0808040001c0400000000000010102000060800080103c12160802000c, sv2v_cast_1(4'h0), 5'h01, 5'h01, 6'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 7'h02, 9'h00c, 7'h04, 10'h020, 7'h07, 5'h01, 10'h027, 8'h08, 9'h004, 8'h0f, 36'h0f0040000, 14'h0004, 6'h02, 7'h03, 5'h01, 7'h05, 9'h001, 6'h02, 8'h01, 5'h01, 5'h01, 7'h01, 7'h03, 6'h03, 8'h08, 7'h02, 8'h05, 8'h03, 5'h01, 18'h00200, 7'h04, 11'h040, 5'h01, 5'h00, 11'h047, 9'h00c, 11'h040, 8'h08, 8'h02, 8'h02, 7'h02, 5'h00, 8'h06, 13'h0010, 7'h01, 5'h01, 17'h00080, 7'h06, 9'h00d, 8'h02, 8'h02, 5'h01, 7'h02, 9'h003, 9'h004, 9'h00c, 5'h01, 5'h00, 8'h08, 9'h004, 5'h01, 8'h0a, 36'h0affff000, 14'h0004, 5'h01, 6'h02, 8'h03, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 36'h000000000, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 5'h00, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 36'h0ffffffff, 5'h00, 5'h00, 5'h01, 6'h02, 8'h03, 9'h004, 7'h02, 9'h00c, 8'h04, 5'h00, 5'h00, 36'h0f00c0000, 9'h00f, 8'h01, 8'h0f, 13'h0020, 12'h01f, 13'h0020, 8'h08, 5'h01, 6'h02, 8'h01, 5'h01};
	input wire [pt[2172-:9]:pt[2163-:6]] hashin;
	input wire [pt[2236-:8] - 1:0] ghr;
	output wire [pt[2270-:8]:pt[2262-:6]] hash;
	generate
		if (pt[2241-:5]) begin : ghrhash_cfg1
			assign hash[pt[2270-:8]:pt[2262-:6]] = {ghr[pt[2236-:8] - 1:pt[2115-:9] - 1], hashin[pt[2115-:9]:2] ^ ghr[pt[2115-:9] - 2:0]};
		end
		else begin : ghrhash_cfg2
			assign hash[pt[2270-:8]:pt[2262-:6]] = {hashin[pt[2236-:8] + 1:2] ^ ghr[pt[2236-:8] - 1:0]};
		end
	endgenerate
endmodule
module rvdff (
	din,
	clk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	output reg [WIDTH - 1:0] dout;
	generate
		if (SHORT == 1) begin
			wire [WIDTH:1] sv2v_tmp_70387;
			assign sv2v_tmp_70387 = din;
			always @(*) dout = sv2v_tmp_70387;
		end
	endgenerate
	always @(posedge clk or negedge rst_l)
		if (rst_l == 0)
			dout[WIDTH - 1:0] <= 0;
		else
			dout[WIDTH - 1:0] <= din[WIDTH - 1:0];
endmodule
module rvdffs (
	din,
	en,
	clk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire en;
	input wire clk;
	input wire rst_l;
	output wire [WIDTH - 1:0] dout;
	generate
		if (SHORT == 1) begin : genblock
			assign dout = din;
		end
		else begin : genblock
			rvdff #(.WIDTH(WIDTH)) dffs(
				.din((en ? din[WIDTH - 1:0] : dout[WIDTH - 1:0])),
				.clk(clk),
				.rst_l(rst_l),
				.dout(dout)
			);
		end
	endgenerate
endmodule
module rvdffsc (
	din,
	en,
	clear,
	clk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire en;
	input wire clear;
	input wire clk;
	input wire rst_l;
	output wire [WIDTH - 1:0] dout;
	wire [WIDTH - 1:0] din_new;
	generate
		if (SHORT == 1) begin
			assign dout = din;
		end
		else begin
			assign din_new = {WIDTH {~clear}} & (en ? din[WIDTH - 1:0] : dout[WIDTH - 1:0]);
			rvdff #(.WIDTH(WIDTH)) dffsc(
				.din(din_new[WIDTH - 1:0]),
				.clk(clk),
				.rst_l(rst_l),
				.dout(dout)
			);
		end
	endgenerate
endmodule
module rvdff_fpga (
	din,
	clk,
	clken,
	rawclk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire clken;
	input wire rawclk;
	input wire rst_l;
	output wire [WIDTH - 1:0] dout;
	generate
		if (SHORT == 1) begin
			assign dout = din;
		end
		else rvdff #(.WIDTH(WIDTH)) dff(
			.din(din),
			.clk(clk),
			.rst_l(rst_l),
			.dout(dout)
		);
	endgenerate
endmodule
module rvdffs_fpga (
	din,
	en,
	clk,
	clken,
	rawclk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire en;
	input wire clk;
	input wire clken;
	input wire rawclk;
	input wire rst_l;
	output wire [WIDTH - 1:0] dout;
	generate
		if (SHORT == 1) begin : genblock
			assign dout = din;
		end
		else begin : genblock
			rvdffs #(.WIDTH(WIDTH)) dffs(
				.din(din),
				.en(en),
				.clk(clk),
				.rst_l(rst_l),
				.dout(dout)
			);
		end
	endgenerate
endmodule
module rvdffsc_fpga (
	din,
	en,
	clear,
	clk,
	clken,
	rawclk,
	rst_l,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	input wire [WIDTH - 1:0] din;
	input wire en;
	input wire clear;
	input wire clk;
	input wire clken;
	input wire rawclk;
	input wire rst_l;
	output wire [WIDTH - 1:0] dout;
	wire [WIDTH - 1:0] din_new;
	generate
		if (SHORT == 1) begin
			assign dout = din;
		end
		else rvdffsc #(.WIDTH(WIDTH)) dffsc(
			.din(din),
			.en(en),
			.clear(clear),
			.clk(clk),
			.rst_l(rst_l),
			.dout(dout)
		);
	endgenerate
endmodule
module rvdffe (
	din,
	en,
	clk,
	rst_l,
	scan_mode,
	dout
);
	parameter WIDTH = 1;
	parameter SHORT = 0;
	parameter OVERRIDE = 0;
	input wire [WIDTH - 1:0] din;
	input wire en;
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	output wire [WIDTH - 1:0] dout;
	wire l1clk;
	generate
		if (SHORT == 1) begin : genblock
			begin : genblock
				assign dout = din;
			end
		end
		else begin : genblock
			rvclkhdr clkhdr(
				.en(en),
				.clk(clk),
				.scan_mode(scan_mode),
				.l1clk(l1clk)
			);
			rvdff #(.WIDTH(WIDTH)) dff(
				.din(din),
				.rst_l(rst_l),
				.dout(dout),
				.clk(l1clk)
			);
		end
	endgenerate
endmodule
module rvdffpcie (
	din,
	clk,
	rst_l,
	en,
	scan_mode,
	dout
);
	parameter WIDTH = 31;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	input wire en;
	input wire scan_mode;
	output wire [WIDTH - 1:0] dout;
	rvdfflie #(
		.WIDTH(WIDTH),
		.LEFT(19)
	) dff(
		.din(din),
		.clk(clk),
		.rst_l(rst_l),
		.en(en),
		.scan_mode(scan_mode),
		.dout(dout)
	);
endmodule
module rvdfflie (
	din,
	clk,
	rst_l,
	en,
	scan_mode,
	dout
);
	parameter WIDTH = 16;
	parameter LEFT = 8;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	input wire en;
	input wire scan_mode;
	output wire [WIDTH - 1:0] dout;
	localparam EXTRA = WIDTH - LEFT;
	localparam LMSB = WIDTH - 1;
	localparam LLSB = (LMSB - LEFT) + 1;
	localparam XMSB = LLSB - 1;
	localparam XLSB = LLSB - EXTRA;
	rvdffiee #(.WIDTH(LEFT)) dff_left(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.en(en),
		.din(din[LMSB:LLSB]),
		.dout(dout[LMSB:LLSB])
	);
	rvdffe #(.WIDTH(EXTRA)) dff_extra(
		.en(en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(din[XMSB:XLSB]),
		.dout(dout[XMSB:XLSB])
	);
endmodule
module rvdffppe (
	din,
	clk,
	rst_l,
	en,
	scan_mode,
	dout
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	input wire en;
	input wire scan_mode;
	output wire [WIDTH - 1:0] dout;
	localparam RIGHT = 31;
	localparam LEFT = WIDTH - RIGHT;
	localparam LMSB = WIDTH - 1;
	localparam LLSB = (LMSB - LEFT) + 1;
	localparam RMSB = LLSB - 1;
	localparam RLSB = LLSB - RIGHT;
	rvdffe #(.WIDTH(LEFT)) dff_left(
		.en(en),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(din[LMSB:LLSB]),
		.dout(dout[LMSB:LLSB])
	);
	rvdffe #(.WIDTH(RIGHT)) dff_right(
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.din(din[RMSB:RLSB]),
		.dout(dout[RMSB:RLSB]),
		.en(en & din[LLSB])
	);
endmodule
module rvdffie (
	din,
	clk,
	rst_l,
	scan_mode,
	dout
);
	parameter WIDTH = 1;
	parameter OVERRIDE = 0;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	output wire [WIDTH - 1:0] dout;
	wire l1clk;
	wire en;
	assign en = |(din ^ dout);
	rvclkhdr clkhdr(
		.en(en),
		.clk(clk),
		.scan_mode(scan_mode),
		.l1clk(l1clk)
	);
	rvdff #(.WIDTH(WIDTH)) dff(
		.din(din),
		.rst_l(rst_l),
		.dout(dout),
		.clk(l1clk)
	);
endmodule
module rvdffiee (
	din,
	clk,
	rst_l,
	scan_mode,
	en,
	dout
);
	parameter WIDTH = 1;
	parameter OVERRIDE = 0;
	input wire [WIDTH - 1:0] din;
	input wire clk;
	input wire rst_l;
	input wire scan_mode;
	input wire en;
	output wire [WIDTH - 1:0] dout;
	wire l1clk;
	wire final_en;
	assign final_en = |(din ^ dout) & en;
	rvdffe #(.WIDTH(WIDTH)) dff(
		.din(din),
		.clk(clk),
		.rst_l(rst_l),
		.scan_mode(scan_mode),
		.dout(dout),
		.en(final_en)
	);
endmodule
module rvsyncss (
	clk,
	rst_l,
	din,
	dout
);
	parameter WIDTH = 251;
	input wire clk;
	input wire rst_l;
	input wire [WIDTH - 1:0] din;
	output wire [WIDTH - 1:0] dout;
	wire [WIDTH - 1:0] din_ff1;
	rvdff #(.WIDTH(WIDTH)) sync_ff1(
		.clk(clk),
		.rst_l(rst_l),
		.din(din[WIDTH - 1:0]),
		.dout(din_ff1[WIDTH - 1:0])
	);
	rvdff #(.WIDTH(WIDTH)) sync_ff2(
		.clk(clk),
		.rst_l(rst_l),
		.din(din_ff1[WIDTH - 1:0]),
		.dout(dout[WIDTH - 1:0])
	);
endmodule
module rvsyncss_fpga (
	gw_clk,
	rawclk,
	clken,
	rst_l,
	din,
	dout
);
	parameter WIDTH = 251;
	input wire gw_clk;
	input wire rawclk;
	input wire clken;
	input wire rst_l;
	input wire [WIDTH - 1:0] din;
	output wire [WIDTH - 1:0] dout;
	wire [WIDTH - 1:0] din_ff1;
	rvdff_fpga #(.WIDTH(WIDTH)) sync_ff1(
		.rst_l(rst_l),
		.clk(gw_clk),
		.rawclk(rawclk),
		.clken(clken),
		.din(din[WIDTH - 1:0]),
		.dout(din_ff1[WIDTH - 1:0])
	);
	rvdff_fpga #(.WIDTH(WIDTH)) sync_ff2(
		.rst_l(rst_l),
		.clk(gw_clk),
		.rawclk(rawclk),
		.clken(clken),
		.din(din_ff1[WIDTH - 1:0]),
		.dout(dout[WIDTH - 1:0])
	);
endmodule
module rvlsadder (
	rs1,
	offset,
	dout
);
	input wire [31:0] rs1;
	input wire [11:0] offset;
	output wire [31:0] dout;
	wire cout;
	wire sign;
	wire [31:12] rs1_inc;
	wire [31:12] rs1_dec;
	assign {cout, dout[11:0]} = {1'b0, rs1[11:0]} + {1'b0, offset[11:0]};
	assign rs1_inc[31:12] = rs1[31:12] + 1;
	assign rs1_dec[31:12] = rs1[31:12] - 1;
	assign sign = offset[11];
	assign dout[31:12] = (({20 {sign ~^ cout}} & rs1[31:12]) | ({20 {~sign & cout}} & rs1_inc[31:12])) | ({20 {sign & ~cout}} & rs1_dec[31:12]);
endmodule
module rvbradder (
	pc,
	offset,
	dout
);
	input [31:1] pc;
	input [12:1] offset;
	output [31:1] dout;
	wire cout;
	wire sign;
	wire [31:13] pc_inc;
	wire [31:13] pc_dec;
	assign {cout, dout[12:1]} = {1'b0, pc[12:1]} + {1'b0, offset[12:1]};
	assign pc_inc[31:13] = pc[31:13] + 1;
	assign pc_dec[31:13] = pc[31:13] - 1;
	assign sign = offset[12];
	assign dout[31:13] = (({19 {sign ~^ cout}} & pc[31:13]) | ({19 {~sign & cout}} & pc_inc[31:13])) | ({19 {sign & ~cout}} & pc_dec[31:13]);
endmodule
module rvtwoscomp (
	din,
	dout
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] din;
	output wire [WIDTH - 1:0] dout;
	wire [WIDTH - 1:1] dout_temp;
	genvar i;
	generate
		for (i = 1; i < WIDTH; i = i + 1) begin : flip_after_first_one
			assign dout_temp[i] = (|din[i - 1:0] ? ~din[i] : din[i]);
		end
	endgenerate
	assign dout[WIDTH - 1:0] = {dout_temp[WIDTH - 1:1], din[0]};
endmodule
module rvfindfirst1 (
	din,
	dout
);
	parameter WIDTH = 32;
	parameter SHIFT = $clog2(WIDTH);
	input wire [WIDTH - 1:0] din;
	output reg [SHIFT - 1:0] dout;
	reg done;
	always @(*) begin
		dout[SHIFT - 1:0] = {SHIFT {1'b0}};
		done = 1'b0;
		begin : sv2v_autoblock_64
			reg signed [31:0] i;
			for (i = WIDTH - 1; i > 0; i = i - 1)
				begin : find_first_one
					done = done | din[i];
					dout[SHIFT - 1:0] = dout[SHIFT - 1:0] + (done ? 1'b0 : 1'b1);
				end
		end
	end
endmodule
module rvfindfirst1hot (
	din,
	dout
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] din;
	output reg [WIDTH - 1:0] dout;
	reg done;
	always @(*) begin
		dout[WIDTH - 1:0] = {WIDTH {1'b0}};
		done = 1'b0;
		begin : sv2v_autoblock_65
			reg signed [31:0] i;
			for (i = 0; i < WIDTH; i = i + 1)
				begin : find_first_one
					dout[i] = ~done & din[i];
					done = done | din[i];
				end
		end
	end
endmodule
module rvmaskandmatch (
	mask,
	data,
	masken,
	match
);
	parameter WIDTH = 32;
	input wire [WIDTH - 1:0] mask;
	input wire [WIDTH - 1:0] data;
	input wire masken;
	output wire match;
	wire [WIDTH - 1:0] matchvec;
	wire masken_or_fullmask;
	assign masken_or_fullmask = masken & ~(&mask[WIDTH - 1:0]);
	assign matchvec[0] = masken_or_fullmask | (mask[0] == data[0]);
	genvar i;
	generate
		for (i = 1; i < WIDTH; i = i + 1) begin : match_after_first_zero
			assign matchvec[i] = (&mask[i - 1:0] & masken_or_fullmask ? 1'b1 : mask[i] == data[i]);
		end
	endgenerate
	assign match = &matchvec[WIDTH - 1:0];
endmodule
module rvrangecheck (
	addr,
	in_range,
	in_region
);
	parameter CCM_SADR = 32'h00000000;
	parameter CCM_SIZE = 128;
	input wire [31:0] addr;
	output wire in_range;
	output wire in_region;
	localparam REGION_BITS = 4;
	localparam MASK_BITS = 10 + $clog2(CCM_SIZE);
	wire [31:0] start_addr;
	wire [3:0] region;
	assign start_addr[31:0] = CCM_SADR;
	assign region[3:0] = start_addr[31:28];
	assign in_region = addr[31:28] == region[3:0];
	generate
		if (CCM_SIZE == 48) begin
			assign in_range = (addr[31:MASK_BITS] == start_addr[31:MASK_BITS]) & ~(&addr[MASK_BITS - 1:MASK_BITS - 2]);
		end
		else assign in_range = addr[31:MASK_BITS] == start_addr[31:MASK_BITS];
	endgenerate
endmodule
module rveven_paritygen (
	data_in,
	parity_out
);
	parameter WIDTH = 16;
	input wire [WIDTH - 1:0] data_in;
	output wire parity_out;
	assign parity_out = ^data_in[WIDTH - 1:0];
endmodule
module rveven_paritycheck (
	data_in,
	parity_in,
	parity_err
);
	parameter WIDTH = 16;
	input wire [WIDTH - 1:0] data_in;
	input wire parity_in;
	output wire parity_err;
	assign parity_err = ^data_in[WIDTH - 1:0] ^ parity_in;
endmodule
module rvecc_encode (
	din,
	ecc_out
);
	input [31:0] din;
	output [6:0] ecc_out;
	wire [5:0] ecc_out_temp;
	assign ecc_out_temp[0] = ((((((((((((((((din[0] ^ din[1]) ^ din[3]) ^ din[4]) ^ din[6]) ^ din[8]) ^ din[10]) ^ din[11]) ^ din[13]) ^ din[15]) ^ din[17]) ^ din[19]) ^ din[21]) ^ din[23]) ^ din[25]) ^ din[26]) ^ din[28]) ^ din[30];
	assign ecc_out_temp[1] = ((((((((((((((((din[0] ^ din[2]) ^ din[3]) ^ din[5]) ^ din[6]) ^ din[9]) ^ din[10]) ^ din[12]) ^ din[13]) ^ din[16]) ^ din[17]) ^ din[20]) ^ din[21]) ^ din[24]) ^ din[25]) ^ din[27]) ^ din[28]) ^ din[31];
	assign ecc_out_temp[2] = ((((((((((((((((din[1] ^ din[2]) ^ din[3]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[29]) ^ din[30]) ^ din[31];
	assign ecc_out_temp[3] = (((((((((((((din[4] ^ din[5]) ^ din[6]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25];
	assign ecc_out_temp[4] = (((((((((((((din[11] ^ din[12]) ^ din[13]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25];
	assign ecc_out_temp[5] = ((((din[26] ^ din[27]) ^ din[28]) ^ din[29]) ^ din[30]) ^ din[31];
	assign ecc_out[6:0] = {^din[31:0] ^ ^ecc_out_temp[5:0], ecc_out_temp[5:0]};
endmodule
module rvecc_decode (
	en,
	din,
	ecc_in,
	sed_ded,
	dout,
	ecc_out,
	single_ecc_error,
	double_ecc_error
);
	input en;
	input [31:0] din;
	input [6:0] ecc_in;
	input sed_ded;
	output [31:0] dout;
	output [6:0] ecc_out;
	output single_ecc_error;
	output double_ecc_error;
	wire [6:0] ecc_check;
	wire [38:0] error_mask;
	wire [38:0] din_plus_parity;
	wire [38:0] dout_plus_parity;
	assign ecc_check[0] = (((((((((((((((((ecc_in[0] ^ din[0]) ^ din[1]) ^ din[3]) ^ din[4]) ^ din[6]) ^ din[8]) ^ din[10]) ^ din[11]) ^ din[13]) ^ din[15]) ^ din[17]) ^ din[19]) ^ din[21]) ^ din[23]) ^ din[25]) ^ din[26]) ^ din[28]) ^ din[30];
	assign ecc_check[1] = (((((((((((((((((ecc_in[1] ^ din[0]) ^ din[2]) ^ din[3]) ^ din[5]) ^ din[6]) ^ din[9]) ^ din[10]) ^ din[12]) ^ din[13]) ^ din[16]) ^ din[17]) ^ din[20]) ^ din[21]) ^ din[24]) ^ din[25]) ^ din[27]) ^ din[28]) ^ din[31];
	assign ecc_check[2] = (((((((((((((((((ecc_in[2] ^ din[1]) ^ din[2]) ^ din[3]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[29]) ^ din[30]) ^ din[31];
	assign ecc_check[3] = ((((((((((((((ecc_in[3] ^ din[4]) ^ din[5]) ^ din[6]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25];
	assign ecc_check[4] = ((((((((((((((ecc_in[4] ^ din[11]) ^ din[12]) ^ din[13]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25];
	assign ecc_check[5] = (((((ecc_in[5] ^ din[26]) ^ din[27]) ^ din[28]) ^ din[29]) ^ din[30]) ^ din[31];
	assign ecc_check[6] = (^din[31:0] ^ ^ecc_in[6:0]) & ~sed_ded;
	assign single_ecc_error = (en & (ecc_check[6:0] != 0)) & ecc_check[6];
	assign double_ecc_error = (en & (ecc_check[6:0] != 0)) & ~ecc_check[6];
	generate
		genvar i;
		for (i = 1; i < 40; i = i + 1) assign error_mask[i - 1] = ecc_check[5:0] == i;
	endgenerate
	assign din_plus_parity[38:0] = {ecc_in[6], din[31:26], ecc_in[5], din[25:11], ecc_in[4], din[10:4], ecc_in[3], din[3:1], ecc_in[2], din[0], ecc_in[1:0]};
	assign dout_plus_parity[38:0] = (single_ecc_error ? error_mask[38:0] ^ din_plus_parity[38:0] : din_plus_parity[38:0]);
	assign dout[31:0] = {dout_plus_parity[37:32], dout_plus_parity[30:16], dout_plus_parity[14:8], dout_plus_parity[6:4], dout_plus_parity[2]};
	assign ecc_out[6:0] = {dout_plus_parity[38] ^ (ecc_check[6:0] == 7'b1000000), dout_plus_parity[31], dout_plus_parity[15], dout_plus_parity[7], dout_plus_parity[3], dout_plus_parity[1:0]};
endmodule
module rvecc_encode_64 (
	din,
	ecc_out
);
	input [63:0] din;
	output [6:0] ecc_out;
	assign ecc_out[0] = (((((((((((((((((((((((((((((((((din[0] ^ din[1]) ^ din[3]) ^ din[4]) ^ din[6]) ^ din[8]) ^ din[10]) ^ din[11]) ^ din[13]) ^ din[15]) ^ din[17]) ^ din[19]) ^ din[21]) ^ din[23]) ^ din[25]) ^ din[26]) ^ din[28]) ^ din[30]) ^ din[32]) ^ din[34]) ^ din[36]) ^ din[38]) ^ din[40]) ^ din[42]) ^ din[44]) ^ din[46]) ^ din[48]) ^ din[50]) ^ din[52]) ^ din[54]) ^ din[56]) ^ din[57]) ^ din[59]) ^ din[61]) ^ din[63];
	assign ecc_out[1] = (((((((((((((((((((((((((((((((((din[0] ^ din[2]) ^ din[3]) ^ din[5]) ^ din[6]) ^ din[9]) ^ din[10]) ^ din[12]) ^ din[13]) ^ din[16]) ^ din[17]) ^ din[20]) ^ din[21]) ^ din[24]) ^ din[25]) ^ din[27]) ^ din[28]) ^ din[31]) ^ din[32]) ^ din[35]) ^ din[36]) ^ din[39]) ^ din[40]) ^ din[43]) ^ din[44]) ^ din[47]) ^ din[48]) ^ din[51]) ^ din[52]) ^ din[55]) ^ din[56]) ^ din[58]) ^ din[59]) ^ din[62]) ^ din[63];
	assign ecc_out[2] = (((((((((((((((((((((((((((((((((din[1] ^ din[2]) ^ din[3]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[29]) ^ din[30]) ^ din[31]) ^ din[32]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56]) ^ din[60]) ^ din[61]) ^ din[62]) ^ din[63];
	assign ecc_out[3] = (((((((((((((((((((((((((((((din[4] ^ din[5]) ^ din[6]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[33]) ^ din[34]) ^ din[35]) ^ din[36]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_out[4] = (((((((((((((((((((((((((((((din[11] ^ din[12]) ^ din[13]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[41]) ^ din[42]) ^ din[43]) ^ din[44]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_out[5] = (((((((((((((((((((((((((((((din[26] ^ din[27]) ^ din[28]) ^ din[29]) ^ din[30]) ^ din[31]) ^ din[32]) ^ din[33]) ^ din[34]) ^ din[35]) ^ din[36]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[41]) ^ din[42]) ^ din[43]) ^ din[44]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_out[6] = (((((din[57] ^ din[58]) ^ din[59]) ^ din[60]) ^ din[61]) ^ din[62]) ^ din[63];
endmodule
module rvecc_decode_64 (
	en,
	din,
	ecc_in,
	ecc_error
);
	input en;
	input [63:0] din;
	input [6:0] ecc_in;
	output ecc_error;
	wire [6:0] ecc_check;
	assign ecc_check[0] = ((((((((((((((((((((((((((((((((((ecc_in[0] ^ din[0]) ^ din[1]) ^ din[3]) ^ din[4]) ^ din[6]) ^ din[8]) ^ din[10]) ^ din[11]) ^ din[13]) ^ din[15]) ^ din[17]) ^ din[19]) ^ din[21]) ^ din[23]) ^ din[25]) ^ din[26]) ^ din[28]) ^ din[30]) ^ din[32]) ^ din[34]) ^ din[36]) ^ din[38]) ^ din[40]) ^ din[42]) ^ din[44]) ^ din[46]) ^ din[48]) ^ din[50]) ^ din[52]) ^ din[54]) ^ din[56]) ^ din[57]) ^ din[59]) ^ din[61]) ^ din[63];
	assign ecc_check[1] = ((((((((((((((((((((((((((((((((((ecc_in[1] ^ din[0]) ^ din[2]) ^ din[3]) ^ din[5]) ^ din[6]) ^ din[9]) ^ din[10]) ^ din[12]) ^ din[13]) ^ din[16]) ^ din[17]) ^ din[20]) ^ din[21]) ^ din[24]) ^ din[25]) ^ din[27]) ^ din[28]) ^ din[31]) ^ din[32]) ^ din[35]) ^ din[36]) ^ din[39]) ^ din[40]) ^ din[43]) ^ din[44]) ^ din[47]) ^ din[48]) ^ din[51]) ^ din[52]) ^ din[55]) ^ din[56]) ^ din[58]) ^ din[59]) ^ din[62]) ^ din[63];
	assign ecc_check[2] = ((((((((((((((((((((((((((((((((((ecc_in[2] ^ din[1]) ^ din[2]) ^ din[3]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[29]) ^ din[30]) ^ din[31]) ^ din[32]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56]) ^ din[60]) ^ din[61]) ^ din[62]) ^ din[63];
	assign ecc_check[3] = ((((((((((((((((((((((((((((((ecc_in[3] ^ din[4]) ^ din[5]) ^ din[6]) ^ din[7]) ^ din[8]) ^ din[9]) ^ din[10]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[33]) ^ din[34]) ^ din[35]) ^ din[36]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_check[4] = ((((((((((((((((((((((((((((((ecc_in[4] ^ din[11]) ^ din[12]) ^ din[13]) ^ din[14]) ^ din[15]) ^ din[16]) ^ din[17]) ^ din[18]) ^ din[19]) ^ din[20]) ^ din[21]) ^ din[22]) ^ din[23]) ^ din[24]) ^ din[25]) ^ din[41]) ^ din[42]) ^ din[43]) ^ din[44]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_check[5] = ((((((((((((((((((((((((((((((ecc_in[5] ^ din[26]) ^ din[27]) ^ din[28]) ^ din[29]) ^ din[30]) ^ din[31]) ^ din[32]) ^ din[33]) ^ din[34]) ^ din[35]) ^ din[36]) ^ din[37]) ^ din[38]) ^ din[39]) ^ din[40]) ^ din[41]) ^ din[42]) ^ din[43]) ^ din[44]) ^ din[45]) ^ din[46]) ^ din[47]) ^ din[48]) ^ din[49]) ^ din[50]) ^ din[51]) ^ din[52]) ^ din[53]) ^ din[54]) ^ din[55]) ^ din[56];
	assign ecc_check[6] = ((((((ecc_in[6] ^ din[57]) ^ din[58]) ^ din[59]) ^ din[60]) ^ din[61]) ^ din[62]) ^ din[63];
	assign ecc_error = en & (ecc_check[6:0] != 0);
endmodule
module rvclkhdr (
	en,
	clk,
	scan_mode,
	l1clk
);
	input wire en;
	input wire clk;
	input wire scan_mode;
	output wire l1clk;
	wire SE;
	assign SE = 0;
	sky130_fd_sc_hd__dlclkp_1 clkhdr(
		.VPWR(1'b1),
		.VGND(1'b0),
		.CLK(clk),
		.GCLK(l1clk),
		.GATE(en)
	);
endmodule
module rvoclkhdr (
	en,
	clk,
	scan_mode,
	l1clk
);
	input wire en;
	input wire clk;
	input wire scan_mode;
	output wire l1clk;
	wire SE;
	assign SE = 0;
	sky130_fd_sc_hd__dlclkp_1 clkhdr(
		.VPWR(1'b1),
		.VGND(1'b0),
		.CLK(clk),
		.GCLK(l1clk),
		.GATE(en)
	);
endmodule
