##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Jun 18 18:35:52 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 2220.420000 BY 3019.880000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540000 0.000000 1.680000 0.485000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300000 0.000000 4.440000 0.485000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.980000 0.000000 468.120000 0.485000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.480000 0.000000 157.620000 0.485000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.580000 0.000000 472.720000 0.485000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.380000 0.000000 463.520000 0.485000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.780000 0.000000 458.920000 0.485000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.640000 0.000000 454.780000 0.485000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.040000 0.000000 450.180000 0.485000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.460000 0.000000 301.600000 0.485000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.860000 0.000000 297.000000 0.485000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.260000 0.000000 292.400000 0.485000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.120000 0.000000 288.260000 0.485000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.520000 0.000000 283.660000 0.485000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.920000 0.000000 279.060000 0.485000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.320000 0.000000 274.460000 0.485000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.720000 0.000000 269.860000 0.485000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.580000 0.000000 265.720000 0.485000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.980000 0.000000 261.120000 0.485000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.380000 0.000000 256.520000 0.485000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.780000 0.000000 251.920000 0.485000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.180000 0.000000 247.320000 0.485000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.040000 0.000000 243.180000 0.485000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.440000 0.000000 238.580000 0.485000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.840000 0.000000 233.980000 0.485000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.240000 0.000000 229.380000 0.485000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.640000 0.000000 224.780000 0.485000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.500000 0.000000 220.640000 0.485000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.900000 0.000000 216.040000 0.485000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300000 0.000000 211.440000 0.485000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.700000 0.000000 206.840000 0.485000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.560000 0.000000 202.700000 0.485000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.960000 0.000000 198.100000 0.485000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360000 0.000000 193.500000 0.485000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.760000 0.000000 188.900000 0.485000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160000 0.000000 184.300000 0.485000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.020000 0.000000 180.160000 0.485000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420000 0.000000 175.560000 0.485000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.820000 0.000000 170.960000 0.485000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220000 0.000000 166.360000 0.485000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620000 0.000000 161.760000 0.485000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.880000 0.000000 153.020000 0.485000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.280000 0.000000 148.420000 0.485000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.680000 0.000000 143.820000 0.485000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080000 0.000000 139.220000 0.485000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.940000 0.000000 135.080000 0.485000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.340000 0.000000 130.480000 0.485000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.740000 0.000000 125.880000 0.485000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.140000 0.000000 121.280000 0.485000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.000000 0.000000 117.140000 0.485000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.400000 0.000000 112.540000 0.485000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.800000 0.000000 107.940000 0.485000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200000 0.000000 103.340000 0.485000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600000 0.000000 98.740000 0.485000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460000 0.000000 94.600000 0.485000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860000 0.000000 90.000000 0.485000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260000 0.000000 85.400000 0.485000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660000 0.000000 80.800000 0.485000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060000 0.000000 76.200000 0.485000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.920000 0.000000 72.060000 0.485000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.320000 0.000000 67.460000 0.485000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720000 0.000000 62.860000 0.485000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.120000 0.000000 58.260000 0.485000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520000 0.000000 53.660000 0.485000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.380000 0.000000 49.520000 0.485000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.780000 0.000000 44.920000 0.485000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180000 0.000000 40.320000 0.485000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580000 0.000000 35.720000 0.485000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.440000 0.000000 31.580000 0.485000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.840000 0.000000 26.980000 0.485000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240000 0.000000 22.380000 0.485000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.640000 0.000000 17.780000 0.485000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040000 0.000000 13.180000 0.485000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900000 0.000000 9.040000 0.485000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.440000 0.000000 445.580000 0.485000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.840000 0.000000 440.980000 0.485000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.700000 0.000000 436.840000 0.485000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.100000 0.000000 432.240000 0.485000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.500000 0.000000 427.640000 0.485000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.900000 0.000000 423.040000 0.485000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.300000 0.000000 418.440000 0.485000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.160000 0.000000 414.300000 0.485000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.560000 0.000000 409.700000 0.485000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.960000 0.000000 405.100000 0.485000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.360000 0.000000 400.500000 0.485000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.760000 0.000000 395.900000 0.485000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.620000 0.000000 391.760000 0.485000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.020000 0.000000 387.160000 0.485000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.420000 0.000000 382.560000 0.485000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.820000 0.000000 377.960000 0.485000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.680000 0.000000 373.820000 0.485000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.080000 0.000000 369.220000 0.485000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.480000 0.000000 364.620000 0.485000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.880000 0.000000 360.020000 0.485000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.280000 0.000000 355.420000 0.485000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.140000 0.000000 351.280000 0.485000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.540000 0.000000 346.680000 0.485000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.940000 0.000000 342.080000 0.485000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.340000 0.000000 337.480000 0.485000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.740000 0.000000 332.880000 0.485000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.600000 0.000000 328.740000 0.485000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.000000 0.000000 324.140000 0.485000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.400000 0.000000 319.540000 0.485000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.800000 0.000000 314.940000 0.485000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.200000 0.000000 310.340000 0.485000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.060000 0.000000 306.200000 0.485000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.960000 0.000000 1049.100000 0.485000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.360000 0.000000 1044.500000 0.485000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.760000 0.000000 1039.900000 0.485000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.620000 0.000000 1035.760000 0.485000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.020000 0.000000 1031.160000 0.485000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.420000 0.000000 1026.560000 0.485000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.820000 0.000000 1021.960000 0.485000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.220000 0.000000 1017.360000 0.485000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.080000 0.000000 1013.220000 0.485000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.480000 0.000000 1008.620000 0.485000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.880000 0.000000 1004.020000 0.485000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.280000 0.000000 999.420000 0.485000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.680000 0.000000 994.820000 0.485000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.540000 0.000000 990.680000 0.485000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.940000 0.000000 986.080000 0.485000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.340000 0.000000 981.480000 0.485000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.740000 0.000000 976.880000 0.485000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.140000 0.000000 972.280000 0.485000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.000000 0.000000 968.140000 0.485000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.400000 0.000000 963.540000 0.485000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.800000 0.000000 958.940000 0.485000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.200000 0.000000 954.340000 0.485000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.060000 0.000000 950.200000 0.485000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.460000 0.000000 945.600000 0.485000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.860000 0.000000 941.000000 0.485000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.260000 0.000000 936.400000 0.485000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.660000 0.000000 931.800000 0.485000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.520000 0.000000 927.660000 0.485000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.920000 0.000000 923.060000 0.485000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.320000 0.000000 918.460000 0.485000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.720000 0.000000 913.860000 0.485000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.120000 0.000000 909.260000 0.485000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.980000 0.000000 905.120000 0.485000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.380000 0.000000 900.520000 0.485000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.780000 0.000000 895.920000 0.485000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.180000 0.000000 891.320000 0.485000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.580000 0.000000 886.720000 0.485000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.440000 0.000000 882.580000 0.485000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.840000 0.000000 877.980000 0.485000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.240000 0.000000 873.380000 0.485000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.640000 0.000000 868.780000 0.485000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.500000 0.000000 864.640000 0.485000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.900000 0.000000 860.040000 0.485000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.300000 0.000000 855.440000 0.485000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.700000 0.000000 850.840000 0.485000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.100000 0.000000 846.240000 0.485000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.960000 0.000000 842.100000 0.485000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.360000 0.000000 837.500000 0.485000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.760000 0.000000 832.900000 0.485000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.160000 0.000000 828.300000 0.485000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.560000 0.000000 823.700000 0.485000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.420000 0.000000 819.560000 0.485000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.820000 0.000000 814.960000 0.485000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.220000 0.000000 810.360000 0.485000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.620000 0.000000 805.760000 0.485000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.020000 0.000000 801.160000 0.485000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.880000 0.000000 797.020000 0.485000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.280000 0.000000 792.420000 0.485000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.680000 0.000000 787.820000 0.485000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.080000 0.000000 783.220000 0.485000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.940000 0.000000 779.080000 0.485000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.340000 0.000000 774.480000 0.485000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.740000 0.000000 769.880000 0.485000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.140000 0.000000 765.280000 0.485000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.540000 0.000000 760.680000 0.485000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.400000 0.000000 756.540000 0.485000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.800000 0.000000 751.940000 0.485000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.200000 0.000000 747.340000 0.485000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.600000 0.000000 742.740000 0.485000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.000000 0.000000 738.140000 0.485000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.860000 0.000000 734.000000 0.485000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.260000 0.000000 729.400000 0.485000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.660000 0.000000 724.800000 0.485000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.060000 0.000000 720.200000 0.485000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.460000 0.000000 715.600000 0.485000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.320000 0.000000 711.460000 0.485000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.720000 0.000000 706.860000 0.485000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.120000 0.000000 702.260000 0.485000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.520000 0.000000 697.660000 0.485000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.380000 0.000000 693.520000 0.485000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.780000 0.000000 688.920000 0.485000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.180000 0.000000 684.320000 0.485000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.580000 0.000000 679.720000 0.485000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.980000 0.000000 675.120000 0.485000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.840000 0.000000 670.980000 0.485000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.240000 0.000000 666.380000 0.485000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.640000 0.000000 661.780000 0.485000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.040000 0.000000 657.180000 0.485000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.440000 0.000000 652.580000 0.485000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.300000 0.000000 648.440000 0.485000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.700000 0.000000 643.840000 0.485000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.100000 0.000000 639.240000 0.485000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.500000 0.000000 634.640000 0.485000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.900000 0.000000 630.040000 0.485000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.760000 0.000000 625.900000 0.485000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.160000 0.000000 621.300000 0.485000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.560000 0.000000 616.700000 0.485000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.960000 0.000000 612.100000 0.485000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.820000 0.000000 607.960000 0.485000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.220000 0.000000 603.360000 0.485000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.620000 0.000000 598.760000 0.485000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.020000 0.000000 594.160000 0.485000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.420000 0.000000 589.560000 0.485000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.280000 0.000000 585.420000 0.485000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.680000 0.000000 580.820000 0.485000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.080000 0.000000 576.220000 0.485000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.480000 0.000000 571.620000 0.485000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.880000 0.000000 567.020000 0.485000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.740000 0.000000 562.880000 0.485000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.140000 0.000000 558.280000 0.485000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.540000 0.000000 553.680000 0.485000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.940000 0.000000 549.080000 0.485000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.340000 0.000000 544.480000 0.485000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.200000 0.000000 540.340000 0.485000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.600000 0.000000 535.740000 0.485000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.000000 0.000000 531.140000 0.485000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.400000 0.000000 526.540000 0.485000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.260000 0.000000 522.400000 0.485000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.660000 0.000000 517.800000 0.485000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.060000 0.000000 513.200000 0.485000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.460000 0.000000 508.600000 0.485000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.860000 0.000000 504.000000 0.485000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.720000 0.000000 499.860000 0.485000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.120000 0.000000 495.260000 0.485000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.520000 0.000000 490.660000 0.485000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.920000 0.000000 486.060000 0.485000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.320000 0.000000 481.460000 0.485000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.180000 0.000000 477.320000 0.485000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.340000 0.000000 1625.480000 0.485000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.740000 0.000000 1620.880000 0.485000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.140000 0.000000 1616.280000 0.485000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.000000 0.000000 1612.140000 0.485000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.400000 0.000000 1607.540000 0.485000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.800000 0.000000 1602.940000 0.485000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.200000 0.000000 1598.340000 0.485000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.600000 0.000000 1593.740000 0.485000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.460000 0.000000 1589.600000 0.485000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.860000 0.000000 1585.000000 0.485000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.260000 0.000000 1580.400000 0.485000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.660000 0.000000 1575.800000 0.485000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.060000 0.000000 1571.200000 0.485000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.920000 0.000000 1567.060000 0.485000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.320000 0.000000 1562.460000 0.485000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.720000 0.000000 1557.860000 0.485000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.120000 0.000000 1553.260000 0.485000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.520000 0.000000 1548.660000 0.485000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.380000 0.000000 1544.520000 0.485000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.780000 0.000000 1539.920000 0.485000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.180000 0.000000 1535.320000 0.485000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.580000 0.000000 1530.720000 0.485000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.440000 0.000000 1526.580000 0.485000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.840000 0.000000 1521.980000 0.485000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.240000 0.000000 1517.380000 0.485000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.640000 0.000000 1512.780000 0.485000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.040000 0.000000 1508.180000 0.485000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.900000 0.000000 1504.040000 0.485000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.300000 0.000000 1499.440000 0.485000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.700000 0.000000 1494.840000 0.485000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.100000 0.000000 1490.240000 0.485000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.500000 0.000000 1485.640000 0.485000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.360000 0.000000 1481.500000 0.485000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.760000 0.000000 1476.900000 0.485000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.160000 0.000000 1472.300000 0.485000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.560000 0.000000 1467.700000 0.485000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.960000 0.000000 1463.100000 0.485000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.820000 0.000000 1458.960000 0.485000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.220000 0.000000 1454.360000 0.485000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.620000 0.000000 1449.760000 0.485000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.020000 0.000000 1445.160000 0.485000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.880000 0.000000 1441.020000 0.485000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.280000 0.000000 1436.420000 0.485000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.680000 0.000000 1431.820000 0.485000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.080000 0.000000 1427.220000 0.485000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.480000 0.000000 1422.620000 0.485000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.340000 0.000000 1418.480000 0.485000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.740000 0.000000 1413.880000 0.485000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.140000 0.000000 1409.280000 0.485000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.540000 0.000000 1404.680000 0.485000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.940000 0.000000 1400.080000 0.485000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.800000 0.000000 1395.940000 0.485000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.200000 0.000000 1391.340000 0.485000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.600000 0.000000 1386.740000 0.485000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.000000 0.000000 1382.140000 0.485000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.400000 0.000000 1377.540000 0.485000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.260000 0.000000 1373.400000 0.485000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.660000 0.000000 1368.800000 0.485000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.060000 0.000000 1364.200000 0.485000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.460000 0.000000 1359.600000 0.485000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.320000 0.000000 1355.460000 0.485000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.720000 0.000000 1350.860000 0.485000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.120000 0.000000 1346.260000 0.485000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.520000 0.000000 1341.660000 0.485000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.920000 0.000000 1337.060000 0.485000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.780000 0.000000 1332.920000 0.485000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.180000 0.000000 1328.320000 0.485000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.580000 0.000000 1323.720000 0.485000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.980000 0.000000 1319.120000 0.485000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.380000 0.000000 1314.520000 0.485000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.240000 0.000000 1310.380000 0.485000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.640000 0.000000 1305.780000 0.485000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.040000 0.000000 1301.180000 0.485000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.440000 0.000000 1296.580000 0.485000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.840000 0.000000 1291.980000 0.485000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.700000 0.000000 1287.840000 0.485000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.100000 0.000000 1283.240000 0.485000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.500000 0.000000 1278.640000 0.485000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.900000 0.000000 1274.040000 0.485000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.760000 0.000000 1269.900000 0.485000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.160000 0.000000 1265.300000 0.485000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.560000 0.000000 1260.700000 0.485000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.960000 0.000000 1256.100000 0.485000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.360000 0.000000 1251.500000 0.485000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.220000 0.000000 1247.360000 0.485000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.620000 0.000000 1242.760000 0.485000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.020000 0.000000 1238.160000 0.485000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.420000 0.000000 1233.560000 0.485000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.820000 0.000000 1228.960000 0.485000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.680000 0.000000 1224.820000 0.485000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.080000 0.000000 1220.220000 0.485000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.480000 0.000000 1215.620000 0.485000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.880000 0.000000 1211.020000 0.485000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.280000 0.000000 1206.420000 0.485000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.140000 0.000000 1202.280000 0.485000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.540000 0.000000 1197.680000 0.485000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.940000 0.000000 1193.080000 0.485000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.340000 0.000000 1188.480000 0.485000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.200000 0.000000 1184.340000 0.485000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.600000 0.000000 1179.740000 0.485000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.000000 0.000000 1175.140000 0.485000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.400000 0.000000 1170.540000 0.485000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.800000 0.000000 1165.940000 0.485000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.660000 0.000000 1161.800000 0.485000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.060000 0.000000 1157.200000 0.485000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.460000 0.000000 1152.600000 0.485000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.860000 0.000000 1148.000000 0.485000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.260000 0.000000 1143.400000 0.485000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.120000 0.000000 1139.260000 0.485000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.520000 0.000000 1134.660000 0.485000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.920000 0.000000 1130.060000 0.485000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.320000 0.000000 1125.460000 0.485000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.720000 0.000000 1120.860000 0.485000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.580000 0.000000 1116.720000 0.485000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.980000 0.000000 1112.120000 0.485000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.380000 0.000000 1107.520000 0.485000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.780000 0.000000 1102.920000 0.485000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.640000 0.000000 1098.780000 0.485000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.040000 0.000000 1094.180000 0.485000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.440000 0.000000 1089.580000 0.485000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.840000 0.000000 1084.980000 0.485000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.240000 0.000000 1080.380000 0.485000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.100000 0.000000 1076.240000 0.485000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.500000 0.000000 1071.640000 0.485000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.900000 0.000000 1067.040000 0.485000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.300000 0.000000 1062.440000 0.485000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.700000 0.000000 1057.840000 0.485000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.560000 0.000000 1053.700000 0.485000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.720000 0.000000 2201.860000 0.485000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.120000 0.000000 2197.260000 0.485000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.520000 0.000000 2192.660000 0.485000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.380000 0.000000 2188.520000 0.485000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.780000 0.000000 2183.920000 0.485000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.180000 0.000000 2179.320000 0.485000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.580000 0.000000 2174.720000 0.485000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2169.980000 0.000000 2170.120000 0.485000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.840000 0.000000 2165.980000 0.485000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.240000 0.000000 2161.380000 0.485000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.640000 0.000000 2156.780000 0.485000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.040000 0.000000 2152.180000 0.485000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.440000 0.000000 2147.580000 0.485000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.300000 0.000000 2143.440000 0.485000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.700000 0.000000 2138.840000 0.485000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.100000 0.000000 2134.240000 0.485000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.500000 0.000000 2129.640000 0.485000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.900000 0.000000 2125.040000 0.485000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.760000 0.000000 2120.900000 0.485000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.160000 0.000000 2116.300000 0.485000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.560000 0.000000 2111.700000 0.485000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.960000 0.000000 2107.100000 0.485000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.820000 0.000000 2102.960000 0.485000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.220000 0.000000 2098.360000 0.485000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.620000 0.000000 2093.760000 0.485000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.020000 0.000000 2089.160000 0.485000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.420000 0.000000 2084.560000 0.485000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.280000 0.000000 2080.420000 0.485000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.680000 0.000000 2075.820000 0.485000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.080000 0.000000 2071.220000 0.485000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.480000 0.000000 2066.620000 0.485000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.880000 0.000000 2062.020000 0.485000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.740000 0.000000 2057.880000 0.485000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.140000 0.000000 2053.280000 0.485000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.540000 0.000000 2048.680000 0.485000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.940000 0.000000 2044.080000 0.485000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.340000 0.000000 2039.480000 0.485000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.200000 0.000000 2035.340000 0.485000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.600000 0.000000 2030.740000 0.485000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.000000 0.000000 2026.140000 0.485000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.400000 0.000000 2021.540000 0.485000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.260000 0.000000 2017.400000 0.485000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.660000 0.000000 2012.800000 0.485000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.060000 0.000000 2008.200000 0.485000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.460000 0.000000 2003.600000 0.485000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.860000 0.000000 1999.000000 0.485000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.720000 0.000000 1994.860000 0.485000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.120000 0.000000 1990.260000 0.485000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.520000 0.000000 1985.660000 0.485000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.920000 0.000000 1981.060000 0.485000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.320000 0.000000 1976.460000 0.485000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.180000 0.000000 1972.320000 0.485000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.580000 0.000000 1967.720000 0.485000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.980000 0.000000 1963.120000 0.485000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.380000 0.000000 1958.520000 0.485000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.780000 0.000000 1953.920000 0.485000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.640000 0.000000 1949.780000 0.485000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.040000 0.000000 1945.180000 0.485000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.440000 0.000000 1940.580000 0.485000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.840000 0.000000 1935.980000 0.485000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.700000 0.000000 1931.840000 0.485000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.100000 0.000000 1927.240000 0.485000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.500000 0.000000 1922.640000 0.485000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.900000 0.000000 1918.040000 0.485000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.300000 0.000000 1913.440000 0.485000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.160000 0.000000 1909.300000 0.485000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.560000 0.000000 1904.700000 0.485000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.960000 0.000000 1900.100000 0.485000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.360000 0.000000 1895.500000 0.485000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.760000 0.000000 1890.900000 0.485000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.620000 0.000000 1886.760000 0.485000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.020000 0.000000 1882.160000 0.485000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.420000 0.000000 1877.560000 0.485000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.820000 0.000000 1872.960000 0.485000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.220000 0.000000 1868.360000 0.485000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.080000 0.000000 1864.220000 0.485000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.480000 0.000000 1859.620000 0.485000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.880000 0.000000 1855.020000 0.485000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.280000 0.000000 1850.420000 0.485000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.140000 0.000000 1846.280000 0.485000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.540000 0.000000 1841.680000 0.485000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.940000 0.000000 1837.080000 0.485000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.340000 0.000000 1832.480000 0.485000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.740000 0.000000 1827.880000 0.485000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.600000 0.000000 1823.740000 0.485000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.000000 0.000000 1819.140000 0.485000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.400000 0.000000 1814.540000 0.485000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.800000 0.000000 1809.940000 0.485000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.200000 0.000000 1805.340000 0.485000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.060000 0.000000 1801.200000 0.485000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.460000 0.000000 1796.600000 0.485000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.860000 0.000000 1792.000000 0.485000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.260000 0.000000 1787.400000 0.485000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.120000 0.000000 1783.260000 0.485000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.520000 0.000000 1778.660000 0.485000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.920000 0.000000 1774.060000 0.485000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.320000 0.000000 1769.460000 0.485000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.720000 0.000000 1764.860000 0.485000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.580000 0.000000 1760.720000 0.485000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.980000 0.000000 1756.120000 0.485000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.380000 0.000000 1751.520000 0.485000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.780000 0.000000 1746.920000 0.485000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.180000 0.000000 1742.320000 0.485000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.040000 0.000000 1738.180000 0.485000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.440000 0.000000 1733.580000 0.485000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.840000 0.000000 1728.980000 0.485000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.240000 0.000000 1724.380000 0.485000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.640000 0.000000 1719.780000 0.485000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.500000 0.000000 1715.640000 0.485000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.900000 0.000000 1711.040000 0.485000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.300000 0.000000 1706.440000 0.485000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.700000 0.000000 1701.840000 0.485000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.560000 0.000000 1697.700000 0.485000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.960000 0.000000 1693.100000 0.485000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.360000 0.000000 1688.500000 0.485000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.760000 0.000000 1683.900000 0.485000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.160000 0.000000 1679.300000 0.485000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.020000 0.000000 1675.160000 0.485000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.420000 0.000000 1670.560000 0.485000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.820000 0.000000 1665.960000 0.485000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.220000 0.000000 1661.360000 0.485000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.620000 0.000000 1656.760000 0.485000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.480000 0.000000 1652.620000 0.485000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.880000 0.000000 1648.020000 0.485000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.280000 0.000000 1643.420000 0.485000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.680000 0.000000 1638.820000 0.485000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.080000 0.000000 1634.220000 0.485000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.940000 0.000000 1630.080000 0.485000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 114.190000 0.800000 114.490000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 284.990000 0.800000 285.290000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 455.790000 0.800000 456.090000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 683.930000 0.800000 684.230000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 912.070000 0.800000 912.370000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1139.600000 0.800000 1139.900000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1367.740000 0.800000 1368.040000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1595.270000 0.800000 1595.570000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1823.410000 0.800000 1823.710000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2051.550000 0.800000 2051.850000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2279.080000 0.800000 2279.380000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2507.220000 0.800000 2507.520000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2735.360000 0.800000 2735.660000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2962.890000 0.800000 2963.190000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.120000 3019.395000 127.260000 3019.880000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.580000 3019.395000 380.720000 3019.880000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.500000 3019.395000 634.640000 3019.880000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.420000 3019.395000 888.560000 3019.880000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.880000 3019.395000 1142.020000 3019.880000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.800000 3019.395000 1395.940000 3019.880000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.720000 3019.395000 1649.860000 3019.880000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.180000 3019.395000 1903.320000 3019.880000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.100000 3019.395000 2157.240000 3019.880000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2903.110000 2220.420000 2903.410000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2670.700000 2220.420000 2671.000000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2438.900000 2220.420000 2439.200000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2206.490000 2220.420000 2206.790000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1974.080000 2220.420000 1974.380000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1741.670000 2220.420000 1741.970000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1509.260000 2220.420000 1509.560000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1277.460000 2220.420000 1277.760000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1045.050000 2220.420000 1045.350000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 870.590000 2220.420000 870.890000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 696.740000 2220.420000 697.040000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 522.280000 2220.420000 522.580000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 347.820000 2220.420000 348.120000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 173.970000 2220.420000 174.270000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1.340000 2220.420000 1.640000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.850000 0.800000 57.150000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 228.260000 0.800000 228.560000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 399.060000 0.800000 399.360000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 627.200000 0.800000 627.500000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 854.730000 0.800000 855.030000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1082.870000 0.800000 1083.170000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1310.400000 0.800000 1310.700000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1538.540000 0.800000 1538.840000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1766.680000 0.800000 1766.980000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1994.210000 0.800000 1994.510000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2222.350000 0.800000 2222.650000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2450.490000 0.800000 2450.790000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2678.020000 0.800000 2678.320000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2906.160000 0.800000 2906.460000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.640000 3019.395000 63.780000 3019.880000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.560000 3019.395000 317.700000 3019.880000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.020000 3019.395000 571.160000 3019.880000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.940000 3019.395000 825.080000 3019.880000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.860000 3019.395000 1079.000000 3019.880000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.320000 3019.395000 1332.460000 3019.880000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.240000 3019.395000 1586.380000 3019.880000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.700000 3019.395000 1839.840000 3019.880000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.620000 3019.395000 2093.760000 3019.880000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2961.060000 2220.420000 2961.360000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2729.260000 2220.420000 2729.560000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2496.850000 2220.420000 2497.150000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2264.440000 2220.420000 2264.740000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2032.030000 2220.420000 2032.330000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1799.620000 2220.420000 1799.920000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1567.820000 2220.420000 1568.120000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1335.410000 2220.420000 1335.710000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1103.000000 2220.420000 1103.300000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 928.540000 2220.420000 928.840000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 754.690000 2220.420000 754.990000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 580.230000 2220.420000 580.530000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 405.770000 2220.420000 406.070000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 231.920000 2220.420000 232.220000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 57.460000 2220.420000 57.760000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2.560000 0.800000 2.860000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 170.920000 0.800000 171.220000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 341.720000 0.800000 342.020000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 569.860000 0.800000 570.160000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 798.000000 0.800000 798.300000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1025.530000 0.800000 1025.830000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1253.670000 0.800000 1253.970000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1481.810000 0.800000 1482.110000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1709.340000 0.800000 1709.640000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1937.480000 0.800000 1937.780000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2165.620000 0.800000 2165.920000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2393.150000 0.800000 2393.450000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2621.290000 0.800000 2621.590000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2848.820000 0.800000 2849.120000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000000 3019.395000 2.140000 3019.880000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.080000 3019.395000 254.220000 3019.880000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.540000 3019.395000 507.680000 3019.880000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.460000 3019.395000 761.600000 3019.880000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.380000 3019.395000 1015.520000 3019.880000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.840000 3019.395000 1268.980000 3019.880000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.760000 3019.395000 1522.900000 3019.880000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.680000 3019.395000 1776.820000 3019.880000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.140000 3019.395000 2030.280000 3019.880000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 3014.740000 2220.420000 3015.040000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2787.210000 2220.420000 2787.510000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2554.800000 2220.420000 2555.100000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2322.390000 2220.420000 2322.690000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2089.980000 2220.420000 2090.280000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1858.180000 2220.420000 1858.480000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1625.770000 2220.420000 1626.070000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1393.360000 2220.420000 1393.660000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1160.950000 2220.420000 1161.250000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 987.100000 2220.420000 987.400000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 812.640000 2220.420000 812.940000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 638.180000 2220.420000 638.480000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 464.330000 2220.420000 464.630000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 289.870000 2220.420000 290.170000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 115.410000 2220.420000 115.710000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 513.130000 0.800000 513.430000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 740.660000 0.800000 740.960000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 968.800000 0.800000 969.100000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1196.940000 0.800000 1197.240000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1424.470000 0.800000 1424.770000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1652.610000 0.800000 1652.910000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1880.140000 0.800000 1880.440000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2108.280000 0.800000 2108.580000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2336.420000 0.800000 2336.720000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2563.950000 0.800000 2564.250000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2792.090000 0.800000 2792.390000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 3015.350000 0.800000 3015.650000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600000 3019.395000 190.740000 3019.880000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.060000 3019.395000 444.200000 3019.880000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.980000 3019.395000 698.120000 3019.880000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.900000 3019.395000 952.040000 3019.880000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.360000 3019.395000 1205.500000 3019.880000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.280000 3019.395000 1459.420000 3019.880000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.200000 3019.395000 1713.340000 3019.880000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.660000 3019.395000 1966.800000 3019.880000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.060000 3019.395000 2215.200000 3019.880000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2845.160000 2220.420000 2845.460000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2612.750000 2220.420000 2613.050000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2380.340000 2220.420000 2380.640000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2148.540000 2220.420000 2148.840000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1916.130000 2220.420000 1916.430000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1683.720000 2220.420000 1684.020000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1451.310000 2220.420000 1451.610000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1218.900000 2220.420000 1219.200000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.320000 0.000000 2206.460000 0.485000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.660000 0.000000 2219.800000 0.485000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.060000 0.000000 2215.200000 0.485000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.460000 0.000000 2210.600000 0.485000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.160000 2.030000 4.160000 3017.849000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1652.635000 2550.185000 1654.375000 2944.965000 ;
      LAYER met4 ;
        RECT 1177.315000 2550.185000 1179.055000 2944.965000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2179.275000 2549.165000 2181.015000 2943.945000 ;
      LAYER met4 ;
        RECT 1703.955000 2549.165000 1705.695000 2943.945000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 634.140000 2550.670000 635.880000 2945.450000 ;
      LAYER met4 ;
        RECT 1109.460000 2550.670000 1111.200000 2945.450000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 72.250000 2550.290000 73.990000 2945.070000 ;
      LAYER met4 ;
        RECT 547.570000 2550.290000 549.310000 2945.070000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2161.300000 34.040000 2163.040000 428.820000 ;
      LAYER met4 ;
        RECT 1685.980000 34.040000 1687.720000 428.820000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1635.570000 19.720000 1637.310000 414.500000 ;
      LAYER met4 ;
        RECT 1160.250000 19.720000 1161.990000 414.500000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1108.280000 26.710000 1110.020000 421.490000 ;
      LAYER met4 ;
        RECT 632.960000 26.710000 634.700000 421.490000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 100.215000 33.220000 101.955000 428.000000 ;
      LAYER met4 ;
        RECT 575.535000 33.220000 577.275000 428.000000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.960000 5.830000 7.960000 3014.050000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1180.715000 2553.585000 1182.455000 2941.565000 ;
      LAYER met4 ;
        RECT 1649.235000 2553.585000 1650.975000 2941.565000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1707.355000 2552.565000 1709.095000 2940.545000 ;
      LAYER met4 ;
        RECT 2175.875000 2552.565000 2177.615000 2940.545000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1106.060000 2554.070000 1107.800000 2942.050000 ;
      LAYER met4 ;
        RECT 637.540000 2554.070000 639.280000 2942.050000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 544.170000 2553.690000 545.910000 2941.670000 ;
      LAYER met4 ;
        RECT 75.650000 2553.690000 77.390000 2941.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1689.380000 37.440000 1691.120000 425.420000 ;
      LAYER met4 ;
        RECT 2157.900000 37.440000 2159.640000 425.420000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1163.650000 23.120000 1165.390000 411.100000 ;
      LAYER met4 ;
        RECT 1632.170000 23.120000 1633.910000 411.100000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 636.360000 30.110000 638.100000 418.090000 ;
      LAYER met4 ;
        RECT 1104.880000 30.110000 1106.620000 418.090000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 572.135000 36.620000 573.875000 424.600000 ;
      LAYER met4 ;
        RECT 103.615000 36.620000 105.355000 424.600000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2220.420000 3019.880000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2220.420000 3019.880000 ;
    LAYER met2 ;
      RECT 2215.340000 3019.255000 2220.420000 3019.880000 ;
      RECT 2157.380000 3019.255000 2214.920000 3019.880000 ;
      RECT 2093.900000 3019.255000 2156.960000 3019.880000 ;
      RECT 2030.420000 3019.255000 2093.480000 3019.880000 ;
      RECT 1966.940000 3019.255000 2030.000000 3019.880000 ;
      RECT 1903.460000 3019.255000 1966.520000 3019.880000 ;
      RECT 1839.980000 3019.255000 1903.040000 3019.880000 ;
      RECT 1776.960000 3019.255000 1839.560000 3019.880000 ;
      RECT 1713.480000 3019.255000 1776.540000 3019.880000 ;
      RECT 1650.000000 3019.255000 1713.060000 3019.880000 ;
      RECT 1586.520000 3019.255000 1649.580000 3019.880000 ;
      RECT 1523.040000 3019.255000 1586.100000 3019.880000 ;
      RECT 1459.560000 3019.255000 1522.620000 3019.880000 ;
      RECT 1396.080000 3019.255000 1459.140000 3019.880000 ;
      RECT 1332.600000 3019.255000 1395.660000 3019.880000 ;
      RECT 1269.120000 3019.255000 1332.180000 3019.880000 ;
      RECT 1205.640000 3019.255000 1268.700000 3019.880000 ;
      RECT 1142.160000 3019.255000 1205.220000 3019.880000 ;
      RECT 1079.140000 3019.255000 1141.740000 3019.880000 ;
      RECT 1015.660000 3019.255000 1078.720000 3019.880000 ;
      RECT 952.180000 3019.255000 1015.240000 3019.880000 ;
      RECT 888.700000 3019.255000 951.760000 3019.880000 ;
      RECT 825.220000 3019.255000 888.280000 3019.880000 ;
      RECT 761.740000 3019.255000 824.800000 3019.880000 ;
      RECT 698.260000 3019.255000 761.320000 3019.880000 ;
      RECT 634.780000 3019.255000 697.840000 3019.880000 ;
      RECT 571.300000 3019.255000 634.360000 3019.880000 ;
      RECT 507.820000 3019.255000 570.880000 3019.880000 ;
      RECT 444.340000 3019.255000 507.400000 3019.880000 ;
      RECT 380.860000 3019.255000 443.920000 3019.880000 ;
      RECT 317.840000 3019.255000 380.440000 3019.880000 ;
      RECT 254.360000 3019.255000 317.420000 3019.880000 ;
      RECT 190.880000 3019.255000 253.940000 3019.880000 ;
      RECT 127.400000 3019.255000 190.460000 3019.880000 ;
      RECT 63.920000 3019.255000 126.980000 3019.880000 ;
      RECT 2.280000 3019.255000 63.500000 3019.880000 ;
      RECT 0.000000 3019.255000 1.860000 3019.880000 ;
      RECT 0.000000 0.625000 2220.420000 3019.255000 ;
      RECT 2219.940000 0.000000 2220.420000 0.625000 ;
      RECT 2215.340000 0.000000 2219.520000 0.625000 ;
      RECT 2210.740000 0.000000 2214.920000 0.625000 ;
      RECT 2206.600000 0.000000 2210.320000 0.625000 ;
      RECT 2202.000000 0.000000 2206.180000 0.625000 ;
      RECT 2197.400000 0.000000 2201.580000 0.625000 ;
      RECT 2192.800000 0.000000 2196.980000 0.625000 ;
      RECT 2188.660000 0.000000 2192.380000 0.625000 ;
      RECT 2184.060000 0.000000 2188.240000 0.625000 ;
      RECT 2179.460000 0.000000 2183.640000 0.625000 ;
      RECT 2174.860000 0.000000 2179.040000 0.625000 ;
      RECT 2170.260000 0.000000 2174.440000 0.625000 ;
      RECT 2166.120000 0.000000 2169.840000 0.625000 ;
      RECT 2161.520000 0.000000 2165.700000 0.625000 ;
      RECT 2156.920000 0.000000 2161.100000 0.625000 ;
      RECT 2152.320000 0.000000 2156.500000 0.625000 ;
      RECT 2147.720000 0.000000 2151.900000 0.625000 ;
      RECT 2143.580000 0.000000 2147.300000 0.625000 ;
      RECT 2138.980000 0.000000 2143.160000 0.625000 ;
      RECT 2134.380000 0.000000 2138.560000 0.625000 ;
      RECT 2129.780000 0.000000 2133.960000 0.625000 ;
      RECT 2125.180000 0.000000 2129.360000 0.625000 ;
      RECT 2121.040000 0.000000 2124.760000 0.625000 ;
      RECT 2116.440000 0.000000 2120.620000 0.625000 ;
      RECT 2111.840000 0.000000 2116.020000 0.625000 ;
      RECT 2107.240000 0.000000 2111.420000 0.625000 ;
      RECT 2103.100000 0.000000 2106.820000 0.625000 ;
      RECT 2098.500000 0.000000 2102.680000 0.625000 ;
      RECT 2093.900000 0.000000 2098.080000 0.625000 ;
      RECT 2089.300000 0.000000 2093.480000 0.625000 ;
      RECT 2084.700000 0.000000 2088.880000 0.625000 ;
      RECT 2080.560000 0.000000 2084.280000 0.625000 ;
      RECT 2075.960000 0.000000 2080.140000 0.625000 ;
      RECT 2071.360000 0.000000 2075.540000 0.625000 ;
      RECT 2066.760000 0.000000 2070.940000 0.625000 ;
      RECT 2062.160000 0.000000 2066.340000 0.625000 ;
      RECT 2058.020000 0.000000 2061.740000 0.625000 ;
      RECT 2053.420000 0.000000 2057.600000 0.625000 ;
      RECT 2048.820000 0.000000 2053.000000 0.625000 ;
      RECT 2044.220000 0.000000 2048.400000 0.625000 ;
      RECT 2039.620000 0.000000 2043.800000 0.625000 ;
      RECT 2035.480000 0.000000 2039.200000 0.625000 ;
      RECT 2030.880000 0.000000 2035.060000 0.625000 ;
      RECT 2026.280000 0.000000 2030.460000 0.625000 ;
      RECT 2021.680000 0.000000 2025.860000 0.625000 ;
      RECT 2017.540000 0.000000 2021.260000 0.625000 ;
      RECT 2012.940000 0.000000 2017.120000 0.625000 ;
      RECT 2008.340000 0.000000 2012.520000 0.625000 ;
      RECT 2003.740000 0.000000 2007.920000 0.625000 ;
      RECT 1999.140000 0.000000 2003.320000 0.625000 ;
      RECT 1995.000000 0.000000 1998.720000 0.625000 ;
      RECT 1990.400000 0.000000 1994.580000 0.625000 ;
      RECT 1985.800000 0.000000 1989.980000 0.625000 ;
      RECT 1981.200000 0.000000 1985.380000 0.625000 ;
      RECT 1976.600000 0.000000 1980.780000 0.625000 ;
      RECT 1972.460000 0.000000 1976.180000 0.625000 ;
      RECT 1967.860000 0.000000 1972.040000 0.625000 ;
      RECT 1963.260000 0.000000 1967.440000 0.625000 ;
      RECT 1958.660000 0.000000 1962.840000 0.625000 ;
      RECT 1954.060000 0.000000 1958.240000 0.625000 ;
      RECT 1949.920000 0.000000 1953.640000 0.625000 ;
      RECT 1945.320000 0.000000 1949.500000 0.625000 ;
      RECT 1940.720000 0.000000 1944.900000 0.625000 ;
      RECT 1936.120000 0.000000 1940.300000 0.625000 ;
      RECT 1931.980000 0.000000 1935.700000 0.625000 ;
      RECT 1927.380000 0.000000 1931.560000 0.625000 ;
      RECT 1922.780000 0.000000 1926.960000 0.625000 ;
      RECT 1918.180000 0.000000 1922.360000 0.625000 ;
      RECT 1913.580000 0.000000 1917.760000 0.625000 ;
      RECT 1909.440000 0.000000 1913.160000 0.625000 ;
      RECT 1904.840000 0.000000 1909.020000 0.625000 ;
      RECT 1900.240000 0.000000 1904.420000 0.625000 ;
      RECT 1895.640000 0.000000 1899.820000 0.625000 ;
      RECT 1891.040000 0.000000 1895.220000 0.625000 ;
      RECT 1886.900000 0.000000 1890.620000 0.625000 ;
      RECT 1882.300000 0.000000 1886.480000 0.625000 ;
      RECT 1877.700000 0.000000 1881.880000 0.625000 ;
      RECT 1873.100000 0.000000 1877.280000 0.625000 ;
      RECT 1868.500000 0.000000 1872.680000 0.625000 ;
      RECT 1864.360000 0.000000 1868.080000 0.625000 ;
      RECT 1859.760000 0.000000 1863.940000 0.625000 ;
      RECT 1855.160000 0.000000 1859.340000 0.625000 ;
      RECT 1850.560000 0.000000 1854.740000 0.625000 ;
      RECT 1846.420000 0.000000 1850.140000 0.625000 ;
      RECT 1841.820000 0.000000 1846.000000 0.625000 ;
      RECT 1837.220000 0.000000 1841.400000 0.625000 ;
      RECT 1832.620000 0.000000 1836.800000 0.625000 ;
      RECT 1828.020000 0.000000 1832.200000 0.625000 ;
      RECT 1823.880000 0.000000 1827.600000 0.625000 ;
      RECT 1819.280000 0.000000 1823.460000 0.625000 ;
      RECT 1814.680000 0.000000 1818.860000 0.625000 ;
      RECT 1810.080000 0.000000 1814.260000 0.625000 ;
      RECT 1805.480000 0.000000 1809.660000 0.625000 ;
      RECT 1801.340000 0.000000 1805.060000 0.625000 ;
      RECT 1796.740000 0.000000 1800.920000 0.625000 ;
      RECT 1792.140000 0.000000 1796.320000 0.625000 ;
      RECT 1787.540000 0.000000 1791.720000 0.625000 ;
      RECT 1783.400000 0.000000 1787.120000 0.625000 ;
      RECT 1778.800000 0.000000 1782.980000 0.625000 ;
      RECT 1774.200000 0.000000 1778.380000 0.625000 ;
      RECT 1769.600000 0.000000 1773.780000 0.625000 ;
      RECT 1765.000000 0.000000 1769.180000 0.625000 ;
      RECT 1760.860000 0.000000 1764.580000 0.625000 ;
      RECT 1756.260000 0.000000 1760.440000 0.625000 ;
      RECT 1751.660000 0.000000 1755.840000 0.625000 ;
      RECT 1747.060000 0.000000 1751.240000 0.625000 ;
      RECT 1742.460000 0.000000 1746.640000 0.625000 ;
      RECT 1738.320000 0.000000 1742.040000 0.625000 ;
      RECT 1733.720000 0.000000 1737.900000 0.625000 ;
      RECT 1729.120000 0.000000 1733.300000 0.625000 ;
      RECT 1724.520000 0.000000 1728.700000 0.625000 ;
      RECT 1719.920000 0.000000 1724.100000 0.625000 ;
      RECT 1715.780000 0.000000 1719.500000 0.625000 ;
      RECT 1711.180000 0.000000 1715.360000 0.625000 ;
      RECT 1706.580000 0.000000 1710.760000 0.625000 ;
      RECT 1701.980000 0.000000 1706.160000 0.625000 ;
      RECT 1697.840000 0.000000 1701.560000 0.625000 ;
      RECT 1693.240000 0.000000 1697.420000 0.625000 ;
      RECT 1688.640000 0.000000 1692.820000 0.625000 ;
      RECT 1684.040000 0.000000 1688.220000 0.625000 ;
      RECT 1679.440000 0.000000 1683.620000 0.625000 ;
      RECT 1675.300000 0.000000 1679.020000 0.625000 ;
      RECT 1670.700000 0.000000 1674.880000 0.625000 ;
      RECT 1666.100000 0.000000 1670.280000 0.625000 ;
      RECT 1661.500000 0.000000 1665.680000 0.625000 ;
      RECT 1656.900000 0.000000 1661.080000 0.625000 ;
      RECT 1652.760000 0.000000 1656.480000 0.625000 ;
      RECT 1648.160000 0.000000 1652.340000 0.625000 ;
      RECT 1643.560000 0.000000 1647.740000 0.625000 ;
      RECT 1638.960000 0.000000 1643.140000 0.625000 ;
      RECT 1634.360000 0.000000 1638.540000 0.625000 ;
      RECT 1630.220000 0.000000 1633.940000 0.625000 ;
      RECT 1625.620000 0.000000 1629.800000 0.625000 ;
      RECT 1621.020000 0.000000 1625.200000 0.625000 ;
      RECT 1616.420000 0.000000 1620.600000 0.625000 ;
      RECT 1612.280000 0.000000 1616.000000 0.625000 ;
      RECT 1607.680000 0.000000 1611.860000 0.625000 ;
      RECT 1603.080000 0.000000 1607.260000 0.625000 ;
      RECT 1598.480000 0.000000 1602.660000 0.625000 ;
      RECT 1593.880000 0.000000 1598.060000 0.625000 ;
      RECT 1589.740000 0.000000 1593.460000 0.625000 ;
      RECT 1585.140000 0.000000 1589.320000 0.625000 ;
      RECT 1580.540000 0.000000 1584.720000 0.625000 ;
      RECT 1575.940000 0.000000 1580.120000 0.625000 ;
      RECT 1571.340000 0.000000 1575.520000 0.625000 ;
      RECT 1567.200000 0.000000 1570.920000 0.625000 ;
      RECT 1562.600000 0.000000 1566.780000 0.625000 ;
      RECT 1558.000000 0.000000 1562.180000 0.625000 ;
      RECT 1553.400000 0.000000 1557.580000 0.625000 ;
      RECT 1548.800000 0.000000 1552.980000 0.625000 ;
      RECT 1544.660000 0.000000 1548.380000 0.625000 ;
      RECT 1540.060000 0.000000 1544.240000 0.625000 ;
      RECT 1535.460000 0.000000 1539.640000 0.625000 ;
      RECT 1530.860000 0.000000 1535.040000 0.625000 ;
      RECT 1526.720000 0.000000 1530.440000 0.625000 ;
      RECT 1522.120000 0.000000 1526.300000 0.625000 ;
      RECT 1517.520000 0.000000 1521.700000 0.625000 ;
      RECT 1512.920000 0.000000 1517.100000 0.625000 ;
      RECT 1508.320000 0.000000 1512.500000 0.625000 ;
      RECT 1504.180000 0.000000 1507.900000 0.625000 ;
      RECT 1499.580000 0.000000 1503.760000 0.625000 ;
      RECT 1494.980000 0.000000 1499.160000 0.625000 ;
      RECT 1490.380000 0.000000 1494.560000 0.625000 ;
      RECT 1485.780000 0.000000 1489.960000 0.625000 ;
      RECT 1481.640000 0.000000 1485.360000 0.625000 ;
      RECT 1477.040000 0.000000 1481.220000 0.625000 ;
      RECT 1472.440000 0.000000 1476.620000 0.625000 ;
      RECT 1467.840000 0.000000 1472.020000 0.625000 ;
      RECT 1463.240000 0.000000 1467.420000 0.625000 ;
      RECT 1459.100000 0.000000 1462.820000 0.625000 ;
      RECT 1454.500000 0.000000 1458.680000 0.625000 ;
      RECT 1449.900000 0.000000 1454.080000 0.625000 ;
      RECT 1445.300000 0.000000 1449.480000 0.625000 ;
      RECT 1441.160000 0.000000 1444.880000 0.625000 ;
      RECT 1436.560000 0.000000 1440.740000 0.625000 ;
      RECT 1431.960000 0.000000 1436.140000 0.625000 ;
      RECT 1427.360000 0.000000 1431.540000 0.625000 ;
      RECT 1422.760000 0.000000 1426.940000 0.625000 ;
      RECT 1418.620000 0.000000 1422.340000 0.625000 ;
      RECT 1414.020000 0.000000 1418.200000 0.625000 ;
      RECT 1409.420000 0.000000 1413.600000 0.625000 ;
      RECT 1404.820000 0.000000 1409.000000 0.625000 ;
      RECT 1400.220000 0.000000 1404.400000 0.625000 ;
      RECT 1396.080000 0.000000 1399.800000 0.625000 ;
      RECT 1391.480000 0.000000 1395.660000 0.625000 ;
      RECT 1386.880000 0.000000 1391.060000 0.625000 ;
      RECT 1382.280000 0.000000 1386.460000 0.625000 ;
      RECT 1377.680000 0.000000 1381.860000 0.625000 ;
      RECT 1373.540000 0.000000 1377.260000 0.625000 ;
      RECT 1368.940000 0.000000 1373.120000 0.625000 ;
      RECT 1364.340000 0.000000 1368.520000 0.625000 ;
      RECT 1359.740000 0.000000 1363.920000 0.625000 ;
      RECT 1355.600000 0.000000 1359.320000 0.625000 ;
      RECT 1351.000000 0.000000 1355.180000 0.625000 ;
      RECT 1346.400000 0.000000 1350.580000 0.625000 ;
      RECT 1341.800000 0.000000 1345.980000 0.625000 ;
      RECT 1337.200000 0.000000 1341.380000 0.625000 ;
      RECT 1333.060000 0.000000 1336.780000 0.625000 ;
      RECT 1328.460000 0.000000 1332.640000 0.625000 ;
      RECT 1323.860000 0.000000 1328.040000 0.625000 ;
      RECT 1319.260000 0.000000 1323.440000 0.625000 ;
      RECT 1314.660000 0.000000 1318.840000 0.625000 ;
      RECT 1310.520000 0.000000 1314.240000 0.625000 ;
      RECT 1305.920000 0.000000 1310.100000 0.625000 ;
      RECT 1301.320000 0.000000 1305.500000 0.625000 ;
      RECT 1296.720000 0.000000 1300.900000 0.625000 ;
      RECT 1292.120000 0.000000 1296.300000 0.625000 ;
      RECT 1287.980000 0.000000 1291.700000 0.625000 ;
      RECT 1283.380000 0.000000 1287.560000 0.625000 ;
      RECT 1278.780000 0.000000 1282.960000 0.625000 ;
      RECT 1274.180000 0.000000 1278.360000 0.625000 ;
      RECT 1270.040000 0.000000 1273.760000 0.625000 ;
      RECT 1265.440000 0.000000 1269.620000 0.625000 ;
      RECT 1260.840000 0.000000 1265.020000 0.625000 ;
      RECT 1256.240000 0.000000 1260.420000 0.625000 ;
      RECT 1251.640000 0.000000 1255.820000 0.625000 ;
      RECT 1247.500000 0.000000 1251.220000 0.625000 ;
      RECT 1242.900000 0.000000 1247.080000 0.625000 ;
      RECT 1238.300000 0.000000 1242.480000 0.625000 ;
      RECT 1233.700000 0.000000 1237.880000 0.625000 ;
      RECT 1229.100000 0.000000 1233.280000 0.625000 ;
      RECT 1224.960000 0.000000 1228.680000 0.625000 ;
      RECT 1220.360000 0.000000 1224.540000 0.625000 ;
      RECT 1215.760000 0.000000 1219.940000 0.625000 ;
      RECT 1211.160000 0.000000 1215.340000 0.625000 ;
      RECT 1206.560000 0.000000 1210.740000 0.625000 ;
      RECT 1202.420000 0.000000 1206.140000 0.625000 ;
      RECT 1197.820000 0.000000 1202.000000 0.625000 ;
      RECT 1193.220000 0.000000 1197.400000 0.625000 ;
      RECT 1188.620000 0.000000 1192.800000 0.625000 ;
      RECT 1184.480000 0.000000 1188.200000 0.625000 ;
      RECT 1179.880000 0.000000 1184.060000 0.625000 ;
      RECT 1175.280000 0.000000 1179.460000 0.625000 ;
      RECT 1170.680000 0.000000 1174.860000 0.625000 ;
      RECT 1166.080000 0.000000 1170.260000 0.625000 ;
      RECT 1161.940000 0.000000 1165.660000 0.625000 ;
      RECT 1157.340000 0.000000 1161.520000 0.625000 ;
      RECT 1152.740000 0.000000 1156.920000 0.625000 ;
      RECT 1148.140000 0.000000 1152.320000 0.625000 ;
      RECT 1143.540000 0.000000 1147.720000 0.625000 ;
      RECT 1139.400000 0.000000 1143.120000 0.625000 ;
      RECT 1134.800000 0.000000 1138.980000 0.625000 ;
      RECT 1130.200000 0.000000 1134.380000 0.625000 ;
      RECT 1125.600000 0.000000 1129.780000 0.625000 ;
      RECT 1121.000000 0.000000 1125.180000 0.625000 ;
      RECT 1116.860000 0.000000 1120.580000 0.625000 ;
      RECT 1112.260000 0.000000 1116.440000 0.625000 ;
      RECT 1107.660000 0.000000 1111.840000 0.625000 ;
      RECT 1103.060000 0.000000 1107.240000 0.625000 ;
      RECT 1098.920000 0.000000 1102.640000 0.625000 ;
      RECT 1094.320000 0.000000 1098.500000 0.625000 ;
      RECT 1089.720000 0.000000 1093.900000 0.625000 ;
      RECT 1085.120000 0.000000 1089.300000 0.625000 ;
      RECT 1080.520000 0.000000 1084.700000 0.625000 ;
      RECT 1076.380000 0.000000 1080.100000 0.625000 ;
      RECT 1071.780000 0.000000 1075.960000 0.625000 ;
      RECT 1067.180000 0.000000 1071.360000 0.625000 ;
      RECT 1062.580000 0.000000 1066.760000 0.625000 ;
      RECT 1057.980000 0.000000 1062.160000 0.625000 ;
      RECT 1053.840000 0.000000 1057.560000 0.625000 ;
      RECT 1049.240000 0.000000 1053.420000 0.625000 ;
      RECT 1044.640000 0.000000 1048.820000 0.625000 ;
      RECT 1040.040000 0.000000 1044.220000 0.625000 ;
      RECT 1035.900000 0.000000 1039.620000 0.625000 ;
      RECT 1031.300000 0.000000 1035.480000 0.625000 ;
      RECT 1026.700000 0.000000 1030.880000 0.625000 ;
      RECT 1022.100000 0.000000 1026.280000 0.625000 ;
      RECT 1017.500000 0.000000 1021.680000 0.625000 ;
      RECT 1013.360000 0.000000 1017.080000 0.625000 ;
      RECT 1008.760000 0.000000 1012.940000 0.625000 ;
      RECT 1004.160000 0.000000 1008.340000 0.625000 ;
      RECT 999.560000 0.000000 1003.740000 0.625000 ;
      RECT 994.960000 0.000000 999.140000 0.625000 ;
      RECT 990.820000 0.000000 994.540000 0.625000 ;
      RECT 986.220000 0.000000 990.400000 0.625000 ;
      RECT 981.620000 0.000000 985.800000 0.625000 ;
      RECT 977.020000 0.000000 981.200000 0.625000 ;
      RECT 972.420000 0.000000 976.600000 0.625000 ;
      RECT 968.280000 0.000000 972.000000 0.625000 ;
      RECT 963.680000 0.000000 967.860000 0.625000 ;
      RECT 959.080000 0.000000 963.260000 0.625000 ;
      RECT 954.480000 0.000000 958.660000 0.625000 ;
      RECT 950.340000 0.000000 954.060000 0.625000 ;
      RECT 945.740000 0.000000 949.920000 0.625000 ;
      RECT 941.140000 0.000000 945.320000 0.625000 ;
      RECT 936.540000 0.000000 940.720000 0.625000 ;
      RECT 931.940000 0.000000 936.120000 0.625000 ;
      RECT 927.800000 0.000000 931.520000 0.625000 ;
      RECT 923.200000 0.000000 927.380000 0.625000 ;
      RECT 918.600000 0.000000 922.780000 0.625000 ;
      RECT 914.000000 0.000000 918.180000 0.625000 ;
      RECT 909.400000 0.000000 913.580000 0.625000 ;
      RECT 905.260000 0.000000 908.980000 0.625000 ;
      RECT 900.660000 0.000000 904.840000 0.625000 ;
      RECT 896.060000 0.000000 900.240000 0.625000 ;
      RECT 891.460000 0.000000 895.640000 0.625000 ;
      RECT 886.860000 0.000000 891.040000 0.625000 ;
      RECT 882.720000 0.000000 886.440000 0.625000 ;
      RECT 878.120000 0.000000 882.300000 0.625000 ;
      RECT 873.520000 0.000000 877.700000 0.625000 ;
      RECT 868.920000 0.000000 873.100000 0.625000 ;
      RECT 864.780000 0.000000 868.500000 0.625000 ;
      RECT 860.180000 0.000000 864.360000 0.625000 ;
      RECT 855.580000 0.000000 859.760000 0.625000 ;
      RECT 850.980000 0.000000 855.160000 0.625000 ;
      RECT 846.380000 0.000000 850.560000 0.625000 ;
      RECT 842.240000 0.000000 845.960000 0.625000 ;
      RECT 837.640000 0.000000 841.820000 0.625000 ;
      RECT 833.040000 0.000000 837.220000 0.625000 ;
      RECT 828.440000 0.000000 832.620000 0.625000 ;
      RECT 823.840000 0.000000 828.020000 0.625000 ;
      RECT 819.700000 0.000000 823.420000 0.625000 ;
      RECT 815.100000 0.000000 819.280000 0.625000 ;
      RECT 810.500000 0.000000 814.680000 0.625000 ;
      RECT 805.900000 0.000000 810.080000 0.625000 ;
      RECT 801.300000 0.000000 805.480000 0.625000 ;
      RECT 797.160000 0.000000 800.880000 0.625000 ;
      RECT 792.560000 0.000000 796.740000 0.625000 ;
      RECT 787.960000 0.000000 792.140000 0.625000 ;
      RECT 783.360000 0.000000 787.540000 0.625000 ;
      RECT 779.220000 0.000000 782.940000 0.625000 ;
      RECT 774.620000 0.000000 778.800000 0.625000 ;
      RECT 770.020000 0.000000 774.200000 0.625000 ;
      RECT 765.420000 0.000000 769.600000 0.625000 ;
      RECT 760.820000 0.000000 765.000000 0.625000 ;
      RECT 756.680000 0.000000 760.400000 0.625000 ;
      RECT 752.080000 0.000000 756.260000 0.625000 ;
      RECT 747.480000 0.000000 751.660000 0.625000 ;
      RECT 742.880000 0.000000 747.060000 0.625000 ;
      RECT 738.280000 0.000000 742.460000 0.625000 ;
      RECT 734.140000 0.000000 737.860000 0.625000 ;
      RECT 729.540000 0.000000 733.720000 0.625000 ;
      RECT 724.940000 0.000000 729.120000 0.625000 ;
      RECT 720.340000 0.000000 724.520000 0.625000 ;
      RECT 715.740000 0.000000 719.920000 0.625000 ;
      RECT 711.600000 0.000000 715.320000 0.625000 ;
      RECT 707.000000 0.000000 711.180000 0.625000 ;
      RECT 702.400000 0.000000 706.580000 0.625000 ;
      RECT 697.800000 0.000000 701.980000 0.625000 ;
      RECT 693.660000 0.000000 697.380000 0.625000 ;
      RECT 689.060000 0.000000 693.240000 0.625000 ;
      RECT 684.460000 0.000000 688.640000 0.625000 ;
      RECT 679.860000 0.000000 684.040000 0.625000 ;
      RECT 675.260000 0.000000 679.440000 0.625000 ;
      RECT 671.120000 0.000000 674.840000 0.625000 ;
      RECT 666.520000 0.000000 670.700000 0.625000 ;
      RECT 661.920000 0.000000 666.100000 0.625000 ;
      RECT 657.320000 0.000000 661.500000 0.625000 ;
      RECT 652.720000 0.000000 656.900000 0.625000 ;
      RECT 648.580000 0.000000 652.300000 0.625000 ;
      RECT 643.980000 0.000000 648.160000 0.625000 ;
      RECT 639.380000 0.000000 643.560000 0.625000 ;
      RECT 634.780000 0.000000 638.960000 0.625000 ;
      RECT 630.180000 0.000000 634.360000 0.625000 ;
      RECT 626.040000 0.000000 629.760000 0.625000 ;
      RECT 621.440000 0.000000 625.620000 0.625000 ;
      RECT 616.840000 0.000000 621.020000 0.625000 ;
      RECT 612.240000 0.000000 616.420000 0.625000 ;
      RECT 608.100000 0.000000 611.820000 0.625000 ;
      RECT 603.500000 0.000000 607.680000 0.625000 ;
      RECT 598.900000 0.000000 603.080000 0.625000 ;
      RECT 594.300000 0.000000 598.480000 0.625000 ;
      RECT 589.700000 0.000000 593.880000 0.625000 ;
      RECT 585.560000 0.000000 589.280000 0.625000 ;
      RECT 580.960000 0.000000 585.140000 0.625000 ;
      RECT 576.360000 0.000000 580.540000 0.625000 ;
      RECT 571.760000 0.000000 575.940000 0.625000 ;
      RECT 567.160000 0.000000 571.340000 0.625000 ;
      RECT 563.020000 0.000000 566.740000 0.625000 ;
      RECT 558.420000 0.000000 562.600000 0.625000 ;
      RECT 553.820000 0.000000 558.000000 0.625000 ;
      RECT 549.220000 0.000000 553.400000 0.625000 ;
      RECT 544.620000 0.000000 548.800000 0.625000 ;
      RECT 540.480000 0.000000 544.200000 0.625000 ;
      RECT 535.880000 0.000000 540.060000 0.625000 ;
      RECT 531.280000 0.000000 535.460000 0.625000 ;
      RECT 526.680000 0.000000 530.860000 0.625000 ;
      RECT 522.540000 0.000000 526.260000 0.625000 ;
      RECT 517.940000 0.000000 522.120000 0.625000 ;
      RECT 513.340000 0.000000 517.520000 0.625000 ;
      RECT 508.740000 0.000000 512.920000 0.625000 ;
      RECT 504.140000 0.000000 508.320000 0.625000 ;
      RECT 500.000000 0.000000 503.720000 0.625000 ;
      RECT 495.400000 0.000000 499.580000 0.625000 ;
      RECT 490.800000 0.000000 494.980000 0.625000 ;
      RECT 486.200000 0.000000 490.380000 0.625000 ;
      RECT 481.600000 0.000000 485.780000 0.625000 ;
      RECT 477.460000 0.000000 481.180000 0.625000 ;
      RECT 472.860000 0.000000 477.040000 0.625000 ;
      RECT 468.260000 0.000000 472.440000 0.625000 ;
      RECT 463.660000 0.000000 467.840000 0.625000 ;
      RECT 459.060000 0.000000 463.240000 0.625000 ;
      RECT 454.920000 0.000000 458.640000 0.625000 ;
      RECT 450.320000 0.000000 454.500000 0.625000 ;
      RECT 445.720000 0.000000 449.900000 0.625000 ;
      RECT 441.120000 0.000000 445.300000 0.625000 ;
      RECT 436.980000 0.000000 440.700000 0.625000 ;
      RECT 432.380000 0.000000 436.560000 0.625000 ;
      RECT 427.780000 0.000000 431.960000 0.625000 ;
      RECT 423.180000 0.000000 427.360000 0.625000 ;
      RECT 418.580000 0.000000 422.760000 0.625000 ;
      RECT 414.440000 0.000000 418.160000 0.625000 ;
      RECT 409.840000 0.000000 414.020000 0.625000 ;
      RECT 405.240000 0.000000 409.420000 0.625000 ;
      RECT 400.640000 0.000000 404.820000 0.625000 ;
      RECT 396.040000 0.000000 400.220000 0.625000 ;
      RECT 391.900000 0.000000 395.620000 0.625000 ;
      RECT 387.300000 0.000000 391.480000 0.625000 ;
      RECT 382.700000 0.000000 386.880000 0.625000 ;
      RECT 378.100000 0.000000 382.280000 0.625000 ;
      RECT 373.960000 0.000000 377.680000 0.625000 ;
      RECT 369.360000 0.000000 373.540000 0.625000 ;
      RECT 364.760000 0.000000 368.940000 0.625000 ;
      RECT 360.160000 0.000000 364.340000 0.625000 ;
      RECT 355.560000 0.000000 359.740000 0.625000 ;
      RECT 351.420000 0.000000 355.140000 0.625000 ;
      RECT 346.820000 0.000000 351.000000 0.625000 ;
      RECT 342.220000 0.000000 346.400000 0.625000 ;
      RECT 337.620000 0.000000 341.800000 0.625000 ;
      RECT 333.020000 0.000000 337.200000 0.625000 ;
      RECT 328.880000 0.000000 332.600000 0.625000 ;
      RECT 324.280000 0.000000 328.460000 0.625000 ;
      RECT 319.680000 0.000000 323.860000 0.625000 ;
      RECT 315.080000 0.000000 319.260000 0.625000 ;
      RECT 310.480000 0.000000 314.660000 0.625000 ;
      RECT 306.340000 0.000000 310.060000 0.625000 ;
      RECT 301.740000 0.000000 305.920000 0.625000 ;
      RECT 297.140000 0.000000 301.320000 0.625000 ;
      RECT 292.540000 0.000000 296.720000 0.625000 ;
      RECT 288.400000 0.000000 292.120000 0.625000 ;
      RECT 283.800000 0.000000 287.980000 0.625000 ;
      RECT 279.200000 0.000000 283.380000 0.625000 ;
      RECT 274.600000 0.000000 278.780000 0.625000 ;
      RECT 270.000000 0.000000 274.180000 0.625000 ;
      RECT 265.860000 0.000000 269.580000 0.625000 ;
      RECT 261.260000 0.000000 265.440000 0.625000 ;
      RECT 256.660000 0.000000 260.840000 0.625000 ;
      RECT 252.060000 0.000000 256.240000 0.625000 ;
      RECT 247.460000 0.000000 251.640000 0.625000 ;
      RECT 243.320000 0.000000 247.040000 0.625000 ;
      RECT 238.720000 0.000000 242.900000 0.625000 ;
      RECT 234.120000 0.000000 238.300000 0.625000 ;
      RECT 229.520000 0.000000 233.700000 0.625000 ;
      RECT 224.920000 0.000000 229.100000 0.625000 ;
      RECT 220.780000 0.000000 224.500000 0.625000 ;
      RECT 216.180000 0.000000 220.360000 0.625000 ;
      RECT 211.580000 0.000000 215.760000 0.625000 ;
      RECT 206.980000 0.000000 211.160000 0.625000 ;
      RECT 202.840000 0.000000 206.560000 0.625000 ;
      RECT 198.240000 0.000000 202.420000 0.625000 ;
      RECT 193.640000 0.000000 197.820000 0.625000 ;
      RECT 189.040000 0.000000 193.220000 0.625000 ;
      RECT 184.440000 0.000000 188.620000 0.625000 ;
      RECT 180.300000 0.000000 184.020000 0.625000 ;
      RECT 175.700000 0.000000 179.880000 0.625000 ;
      RECT 171.100000 0.000000 175.280000 0.625000 ;
      RECT 166.500000 0.000000 170.680000 0.625000 ;
      RECT 161.900000 0.000000 166.080000 0.625000 ;
      RECT 157.760000 0.000000 161.480000 0.625000 ;
      RECT 153.160000 0.000000 157.340000 0.625000 ;
      RECT 148.560000 0.000000 152.740000 0.625000 ;
      RECT 143.960000 0.000000 148.140000 0.625000 ;
      RECT 139.360000 0.000000 143.540000 0.625000 ;
      RECT 135.220000 0.000000 138.940000 0.625000 ;
      RECT 130.620000 0.000000 134.800000 0.625000 ;
      RECT 126.020000 0.000000 130.200000 0.625000 ;
      RECT 121.420000 0.000000 125.600000 0.625000 ;
      RECT 117.280000 0.000000 121.000000 0.625000 ;
      RECT 112.680000 0.000000 116.860000 0.625000 ;
      RECT 108.080000 0.000000 112.260000 0.625000 ;
      RECT 103.480000 0.000000 107.660000 0.625000 ;
      RECT 98.880000 0.000000 103.060000 0.625000 ;
      RECT 94.740000 0.000000 98.460000 0.625000 ;
      RECT 90.140000 0.000000 94.320000 0.625000 ;
      RECT 85.540000 0.000000 89.720000 0.625000 ;
      RECT 80.940000 0.000000 85.120000 0.625000 ;
      RECT 76.340000 0.000000 80.520000 0.625000 ;
      RECT 72.200000 0.000000 75.920000 0.625000 ;
      RECT 67.600000 0.000000 71.780000 0.625000 ;
      RECT 63.000000 0.000000 67.180000 0.625000 ;
      RECT 58.400000 0.000000 62.580000 0.625000 ;
      RECT 53.800000 0.000000 57.980000 0.625000 ;
      RECT 49.660000 0.000000 53.380000 0.625000 ;
      RECT 45.060000 0.000000 49.240000 0.625000 ;
      RECT 40.460000 0.000000 44.640000 0.625000 ;
      RECT 35.860000 0.000000 40.040000 0.625000 ;
      RECT 31.720000 0.000000 35.440000 0.625000 ;
      RECT 27.120000 0.000000 31.300000 0.625000 ;
      RECT 22.520000 0.000000 26.700000 0.625000 ;
      RECT 17.920000 0.000000 22.100000 0.625000 ;
      RECT 13.320000 0.000000 17.500000 0.625000 ;
      RECT 9.180000 0.000000 12.900000 0.625000 ;
      RECT 4.580000 0.000000 8.760000 0.625000 ;
      RECT 1.820000 0.000000 4.160000 0.625000 ;
      RECT 0.000000 0.000000 1.400000 0.625000 ;
    LAYER met3 ;
      RECT 0.000000 3015.950000 2220.420000 3019.880000 ;
      RECT 1.100000 3015.340000 2220.420000 3015.950000 ;
      RECT 1.100000 3015.050000 2219.320000 3015.340000 ;
      RECT 0.000000 3014.440000 2219.320000 3015.050000 ;
      RECT 0.000000 2963.490000 2220.420000 3014.440000 ;
      RECT 1.100000 2962.590000 2220.420000 2963.490000 ;
      RECT 0.000000 2961.660000 2220.420000 2962.590000 ;
      RECT 0.000000 2960.760000 2219.320000 2961.660000 ;
      RECT 0.000000 2906.760000 2220.420000 2960.760000 ;
      RECT 1.100000 2905.860000 2220.420000 2906.760000 ;
      RECT 0.000000 2903.710000 2220.420000 2905.860000 ;
      RECT 0.000000 2902.810000 2219.320000 2903.710000 ;
      RECT 0.000000 2849.420000 2220.420000 2902.810000 ;
      RECT 1.100000 2848.520000 2220.420000 2849.420000 ;
      RECT 0.000000 2845.760000 2220.420000 2848.520000 ;
      RECT 0.000000 2844.860000 2219.320000 2845.760000 ;
      RECT 0.000000 2792.690000 2220.420000 2844.860000 ;
      RECT 1.100000 2791.790000 2220.420000 2792.690000 ;
      RECT 0.000000 2787.810000 2220.420000 2791.790000 ;
      RECT 0.000000 2786.910000 2219.320000 2787.810000 ;
      RECT 0.000000 2735.960000 2220.420000 2786.910000 ;
      RECT 1.100000 2735.060000 2220.420000 2735.960000 ;
      RECT 0.000000 2729.860000 2220.420000 2735.060000 ;
      RECT 0.000000 2728.960000 2219.320000 2729.860000 ;
      RECT 0.000000 2678.620000 2220.420000 2728.960000 ;
      RECT 1.100000 2677.720000 2220.420000 2678.620000 ;
      RECT 0.000000 2671.300000 2220.420000 2677.720000 ;
      RECT 0.000000 2670.400000 2219.320000 2671.300000 ;
      RECT 0.000000 2621.890000 2220.420000 2670.400000 ;
      RECT 1.100000 2620.990000 2220.420000 2621.890000 ;
      RECT 0.000000 2613.350000 2220.420000 2620.990000 ;
      RECT 0.000000 2612.450000 2219.320000 2613.350000 ;
      RECT 0.000000 2564.550000 2220.420000 2612.450000 ;
      RECT 1.100000 2563.650000 2220.420000 2564.550000 ;
      RECT 0.000000 2555.400000 2220.420000 2563.650000 ;
      RECT 0.000000 2554.500000 2219.320000 2555.400000 ;
      RECT 0.000000 2507.820000 2220.420000 2554.500000 ;
      RECT 1.100000 2506.920000 2220.420000 2507.820000 ;
      RECT 0.000000 2497.450000 2220.420000 2506.920000 ;
      RECT 0.000000 2496.550000 2219.320000 2497.450000 ;
      RECT 0.000000 2451.090000 2220.420000 2496.550000 ;
      RECT 1.100000 2450.190000 2220.420000 2451.090000 ;
      RECT 0.000000 2439.500000 2220.420000 2450.190000 ;
      RECT 0.000000 2438.600000 2219.320000 2439.500000 ;
      RECT 0.000000 2393.750000 2220.420000 2438.600000 ;
      RECT 1.100000 2392.850000 2220.420000 2393.750000 ;
      RECT 0.000000 2380.940000 2220.420000 2392.850000 ;
      RECT 0.000000 2380.040000 2219.320000 2380.940000 ;
      RECT 0.000000 2337.020000 2220.420000 2380.040000 ;
      RECT 1.100000 2336.120000 2220.420000 2337.020000 ;
      RECT 0.000000 2322.990000 2220.420000 2336.120000 ;
      RECT 0.000000 2322.090000 2219.320000 2322.990000 ;
      RECT 0.000000 2279.680000 2220.420000 2322.090000 ;
      RECT 1.100000 2278.780000 2220.420000 2279.680000 ;
      RECT 0.000000 2265.040000 2220.420000 2278.780000 ;
      RECT 0.000000 2264.140000 2219.320000 2265.040000 ;
      RECT 0.000000 2222.950000 2220.420000 2264.140000 ;
      RECT 1.100000 2222.050000 2220.420000 2222.950000 ;
      RECT 0.000000 2207.090000 2220.420000 2222.050000 ;
      RECT 0.000000 2206.190000 2219.320000 2207.090000 ;
      RECT 0.000000 2166.220000 2220.420000 2206.190000 ;
      RECT 1.100000 2165.320000 2220.420000 2166.220000 ;
      RECT 0.000000 2149.140000 2220.420000 2165.320000 ;
      RECT 0.000000 2148.240000 2219.320000 2149.140000 ;
      RECT 0.000000 2108.880000 2220.420000 2148.240000 ;
      RECT 1.100000 2107.980000 2220.420000 2108.880000 ;
      RECT 0.000000 2090.580000 2220.420000 2107.980000 ;
      RECT 0.000000 2089.680000 2219.320000 2090.580000 ;
      RECT 0.000000 2052.150000 2220.420000 2089.680000 ;
      RECT 1.100000 2051.250000 2220.420000 2052.150000 ;
      RECT 0.000000 2032.630000 2220.420000 2051.250000 ;
      RECT 0.000000 2031.730000 2219.320000 2032.630000 ;
      RECT 0.000000 1994.810000 2220.420000 2031.730000 ;
      RECT 1.100000 1993.910000 2220.420000 1994.810000 ;
      RECT 0.000000 1974.680000 2220.420000 1993.910000 ;
      RECT 0.000000 1973.780000 2219.320000 1974.680000 ;
      RECT 0.000000 1938.080000 2220.420000 1973.780000 ;
      RECT 1.100000 1937.180000 2220.420000 1938.080000 ;
      RECT 0.000000 1916.730000 2220.420000 1937.180000 ;
      RECT 0.000000 1915.830000 2219.320000 1916.730000 ;
      RECT 0.000000 1880.740000 2220.420000 1915.830000 ;
      RECT 1.100000 1879.840000 2220.420000 1880.740000 ;
      RECT 0.000000 1858.780000 2220.420000 1879.840000 ;
      RECT 0.000000 1857.880000 2219.320000 1858.780000 ;
      RECT 0.000000 1824.010000 2220.420000 1857.880000 ;
      RECT 1.100000 1823.110000 2220.420000 1824.010000 ;
      RECT 0.000000 1800.220000 2220.420000 1823.110000 ;
      RECT 0.000000 1799.320000 2219.320000 1800.220000 ;
      RECT 0.000000 1767.280000 2220.420000 1799.320000 ;
      RECT 1.100000 1766.380000 2220.420000 1767.280000 ;
      RECT 0.000000 1742.270000 2220.420000 1766.380000 ;
      RECT 0.000000 1741.370000 2219.320000 1742.270000 ;
      RECT 0.000000 1709.940000 2220.420000 1741.370000 ;
      RECT 1.100000 1709.040000 2220.420000 1709.940000 ;
      RECT 0.000000 1684.320000 2220.420000 1709.040000 ;
      RECT 0.000000 1683.420000 2219.320000 1684.320000 ;
      RECT 0.000000 1653.210000 2220.420000 1683.420000 ;
      RECT 1.100000 1652.310000 2220.420000 1653.210000 ;
      RECT 0.000000 1626.370000 2220.420000 1652.310000 ;
      RECT 0.000000 1625.470000 2219.320000 1626.370000 ;
      RECT 0.000000 1595.870000 2220.420000 1625.470000 ;
      RECT 1.100000 1594.970000 2220.420000 1595.870000 ;
      RECT 0.000000 1568.420000 2220.420000 1594.970000 ;
      RECT 0.000000 1567.520000 2219.320000 1568.420000 ;
      RECT 0.000000 1539.140000 2220.420000 1567.520000 ;
      RECT 1.100000 1538.240000 2220.420000 1539.140000 ;
      RECT 0.000000 1509.860000 2220.420000 1538.240000 ;
      RECT 0.000000 1508.960000 2219.320000 1509.860000 ;
      RECT 0.000000 1482.410000 2220.420000 1508.960000 ;
      RECT 1.100000 1481.510000 2220.420000 1482.410000 ;
      RECT 0.000000 1451.910000 2220.420000 1481.510000 ;
      RECT 0.000000 1451.010000 2219.320000 1451.910000 ;
      RECT 0.000000 1425.070000 2220.420000 1451.010000 ;
      RECT 1.100000 1424.170000 2220.420000 1425.070000 ;
      RECT 0.000000 1393.960000 2220.420000 1424.170000 ;
      RECT 0.000000 1393.060000 2219.320000 1393.960000 ;
      RECT 0.000000 1368.340000 2220.420000 1393.060000 ;
      RECT 1.100000 1367.440000 2220.420000 1368.340000 ;
      RECT 0.000000 1336.010000 2220.420000 1367.440000 ;
      RECT 0.000000 1335.110000 2219.320000 1336.010000 ;
      RECT 0.000000 1311.000000 2220.420000 1335.110000 ;
      RECT 1.100000 1310.100000 2220.420000 1311.000000 ;
      RECT 0.000000 1278.060000 2220.420000 1310.100000 ;
      RECT 0.000000 1277.160000 2219.320000 1278.060000 ;
      RECT 0.000000 1254.270000 2220.420000 1277.160000 ;
      RECT 1.100000 1253.370000 2220.420000 1254.270000 ;
      RECT 0.000000 1219.500000 2220.420000 1253.370000 ;
      RECT 0.000000 1218.600000 2219.320000 1219.500000 ;
      RECT 0.000000 1197.540000 2220.420000 1218.600000 ;
      RECT 1.100000 1196.640000 2220.420000 1197.540000 ;
      RECT 0.000000 1161.550000 2220.420000 1196.640000 ;
      RECT 0.000000 1160.650000 2219.320000 1161.550000 ;
      RECT 0.000000 1140.200000 2220.420000 1160.650000 ;
      RECT 1.100000 1139.300000 2220.420000 1140.200000 ;
      RECT 0.000000 1103.600000 2220.420000 1139.300000 ;
      RECT 0.000000 1102.700000 2219.320000 1103.600000 ;
      RECT 0.000000 1083.470000 2220.420000 1102.700000 ;
      RECT 1.100000 1082.570000 2220.420000 1083.470000 ;
      RECT 0.000000 1045.650000 2220.420000 1082.570000 ;
      RECT 0.000000 1044.750000 2219.320000 1045.650000 ;
      RECT 0.000000 1026.130000 2220.420000 1044.750000 ;
      RECT 1.100000 1025.230000 2220.420000 1026.130000 ;
      RECT 0.000000 987.700000 2220.420000 1025.230000 ;
      RECT 0.000000 986.800000 2219.320000 987.700000 ;
      RECT 0.000000 969.400000 2220.420000 986.800000 ;
      RECT 1.100000 968.500000 2220.420000 969.400000 ;
      RECT 0.000000 929.140000 2220.420000 968.500000 ;
      RECT 0.000000 928.240000 2219.320000 929.140000 ;
      RECT 0.000000 912.670000 2220.420000 928.240000 ;
      RECT 1.100000 911.770000 2220.420000 912.670000 ;
      RECT 0.000000 871.190000 2220.420000 911.770000 ;
      RECT 0.000000 870.290000 2219.320000 871.190000 ;
      RECT 0.000000 855.330000 2220.420000 870.290000 ;
      RECT 1.100000 854.430000 2220.420000 855.330000 ;
      RECT 0.000000 813.240000 2220.420000 854.430000 ;
      RECT 0.000000 812.340000 2219.320000 813.240000 ;
      RECT 0.000000 798.600000 2220.420000 812.340000 ;
      RECT 1.100000 797.700000 2220.420000 798.600000 ;
      RECT 0.000000 755.290000 2220.420000 797.700000 ;
      RECT 0.000000 754.390000 2219.320000 755.290000 ;
      RECT 0.000000 741.260000 2220.420000 754.390000 ;
      RECT 1.100000 740.360000 2220.420000 741.260000 ;
      RECT 0.000000 697.340000 2220.420000 740.360000 ;
      RECT 0.000000 696.440000 2219.320000 697.340000 ;
      RECT 0.000000 684.530000 2220.420000 696.440000 ;
      RECT 1.100000 683.630000 2220.420000 684.530000 ;
      RECT 0.000000 638.780000 2220.420000 683.630000 ;
      RECT 0.000000 637.880000 2219.320000 638.780000 ;
      RECT 0.000000 627.800000 2220.420000 637.880000 ;
      RECT 1.100000 626.900000 2220.420000 627.800000 ;
      RECT 0.000000 580.830000 2220.420000 626.900000 ;
      RECT 0.000000 579.930000 2219.320000 580.830000 ;
      RECT 0.000000 570.460000 2220.420000 579.930000 ;
      RECT 1.100000 569.560000 2220.420000 570.460000 ;
      RECT 0.000000 522.880000 2220.420000 569.560000 ;
      RECT 0.000000 521.980000 2219.320000 522.880000 ;
      RECT 0.000000 513.730000 2220.420000 521.980000 ;
      RECT 1.100000 512.830000 2220.420000 513.730000 ;
      RECT 0.000000 464.930000 2220.420000 512.830000 ;
      RECT 0.000000 464.030000 2219.320000 464.930000 ;
      RECT 0.000000 456.390000 2220.420000 464.030000 ;
      RECT 1.100000 455.490000 2220.420000 456.390000 ;
      RECT 0.000000 406.370000 2220.420000 455.490000 ;
      RECT 0.000000 405.470000 2219.320000 406.370000 ;
      RECT 0.000000 399.660000 2220.420000 405.470000 ;
      RECT 1.100000 398.760000 2220.420000 399.660000 ;
      RECT 0.000000 348.420000 2220.420000 398.760000 ;
      RECT 0.000000 347.520000 2219.320000 348.420000 ;
      RECT 0.000000 342.320000 2220.420000 347.520000 ;
      RECT 1.100000 341.420000 2220.420000 342.320000 ;
      RECT 0.000000 290.470000 2220.420000 341.420000 ;
      RECT 0.000000 289.570000 2219.320000 290.470000 ;
      RECT 0.000000 285.590000 2220.420000 289.570000 ;
      RECT 1.100000 284.690000 2220.420000 285.590000 ;
      RECT 0.000000 232.520000 2220.420000 284.690000 ;
      RECT 0.000000 231.620000 2219.320000 232.520000 ;
      RECT 0.000000 228.860000 2220.420000 231.620000 ;
      RECT 1.100000 227.960000 2220.420000 228.860000 ;
      RECT 0.000000 174.570000 2220.420000 227.960000 ;
      RECT 0.000000 173.670000 2219.320000 174.570000 ;
      RECT 0.000000 171.520000 2220.420000 173.670000 ;
      RECT 1.100000 170.620000 2220.420000 171.520000 ;
      RECT 0.000000 116.010000 2220.420000 170.620000 ;
      RECT 0.000000 115.110000 2219.320000 116.010000 ;
      RECT 0.000000 114.790000 2220.420000 115.110000 ;
      RECT 1.100000 113.890000 2220.420000 114.790000 ;
      RECT 0.000000 58.060000 2220.420000 113.890000 ;
      RECT 0.000000 57.450000 2219.320000 58.060000 ;
      RECT 1.100000 57.160000 2219.320000 57.450000 ;
      RECT 1.100000 56.550000 2220.420000 57.160000 ;
      RECT 0.000000 3.160000 2220.420000 56.550000 ;
      RECT 1.100000 2.260000 2220.420000 3.160000 ;
      RECT 0.000000 1.940000 2220.420000 2.260000 ;
      RECT 0.000000 1.040000 2219.320000 1.940000 ;
      RECT 0.000000 0.000000 2220.420000 1.040000 ;
    LAYER met4 ;
      RECT 0.000000 3018.149000 2220.420000 3019.880000 ;
      RECT 4.460000 3014.350000 2220.420000 3018.149000 ;
      RECT 8.260000 5.530000 2220.420000 3014.350000 ;
      RECT 4.460000 5.530000 5.660000 3014.350000 ;
      RECT 4.460000 1.730000 2220.420000 5.530000 ;
      RECT 0.000000 1.730000 1.860000 3018.149000 ;
      RECT 0.000000 0.000000 2220.420000 1.730000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2220.420000 3019.880000 ;
  END
END user_proj_example

END LIBRARY
