magic
tech sky130A
magscale 1 2
timestamp 1625000815
<< locali >>
rect 292313 11033 292497 11067
rect 292313 10999 292347 11033
rect 302283 10965 302467 10999
rect 277593 10455 277627 10761
rect 282837 10455 282871 10965
rect 286885 10591 286919 10761
rect 286885 10557 287253 10591
rect 287621 10523 287655 10557
rect 292405 10523 292439 10965
rect 302283 10761 302375 10795
rect 287621 10489 287805 10523
rect 292347 10489 292439 10523
rect 277593 10421 278145 10455
rect 282779 10421 282871 10455
rect 302341 10183 302375 10761
rect 302433 10523 302467 10965
rect 306389 10523 306423 10557
rect 306239 10489 306423 10523
rect 302249 9639 302283 10149
rect 306941 10115 306975 10557
rect 307217 10183 307251 10693
rect 311633 10591 311667 10625
rect 311633 10557 311909 10591
rect 311541 10523 311575 10557
rect 311541 10489 311817 10523
rect 307309 10115 307343 10149
rect 306941 10081 307343 10115
rect 307125 9979 307159 10013
rect 306975 9945 307159 9979
rect 284125 9367 284159 9469
rect 292313 9469 292497 9503
rect 284125 9333 284401 9367
rect 287529 9027 287563 9333
rect 287621 9095 287655 9333
rect 292313 9163 292347 9469
rect 292405 9129 292497 9163
rect 292405 9027 292439 9129
rect 287529 8993 287805 9027
rect 253213 8075 253247 8245
rect 253305 7735 253339 8041
rect 253489 7395 253523 7769
rect 292497 7395 292531 8993
rect 400045 7191 400079 7293
rect 400045 7157 400321 7191
rect 348927 6681 349387 6715
rect 349353 6443 349387 6681
rect 398113 6647 398147 6749
rect 394525 6443 394559 6613
rect 398021 6579 398055 6613
rect 398205 6579 398239 6749
rect 398021 6545 398239 6579
rect 394433 6307 394467 6409
rect 394433 6273 394801 6307
rect 209421 5287 209455 5593
rect 209513 5219 209547 5525
rect 209605 5151 209639 5253
rect 209421 5117 209639 5151
rect 209421 4811 209455 5117
rect 209697 5015 209731 5185
rect 219633 5083 219667 5593
rect 219725 5151 219759 5525
rect 277041 5355 277075 5593
rect 320741 5559 320775 5661
rect 327733 5559 327767 5797
rect 349905 5627 349939 6273
rect 463893 6239 463927 7497
rect 465733 6919 465767 7361
rect 465825 6919 465859 7497
rect 278271 5253 278421 5287
rect 279709 5219 279743 5525
rect 282653 5355 282687 5525
rect 320833 5525 321017 5559
rect 388453 5559 388487 6205
rect 463709 6171 463743 6205
rect 463985 6171 464019 6205
rect 463709 6137 464019 6171
rect 502257 6171 502291 6885
rect 320649 5491 320683 5525
rect 320833 5491 320867 5525
rect 320649 5457 320867 5491
rect 209547 4981 209731 5015
rect 34529 3383 34563 3553
rect 92489 3179 92523 3349
rect 116317 2839 116351 3689
rect 123217 2839 123251 4165
rect 124597 3519 124631 3689
rect 128553 3655 128587 4165
rect 123309 2839 123343 3417
rect 126897 2635 126931 3485
rect 127633 3451 127667 3621
rect 127541 3383 127575 3417
rect 127725 3383 127759 3621
rect 132785 3519 132819 4165
rect 219541 4131 219575 5049
rect 277903 4709 278087 4743
rect 278053 4675 278087 4709
rect 278145 4607 278179 5185
rect 509341 5015 509375 5525
rect 132877 3519 132911 4029
rect 451323 3893 451415 3927
rect 451381 3723 451415 3893
rect 455429 3723 455463 3893
rect 128461 3451 128495 3485
rect 128461 3417 128645 3451
rect 127541 3349 127759 3383
rect 156981 3383 157015 3485
rect 158579 3417 158729 3451
rect 426081 2975 426115 3621
rect 128461 2567 128495 2805
rect 436695 2805 437489 2839
rect 132325 2635 132359 2805
rect 460765 2635 460799 3893
rect 461041 3383 461075 4029
rect 460949 3111 460983 3349
rect 460949 3077 461225 3111
rect 461317 3043 461351 4097
rect 461501 4029 462513 4063
rect 461501 3451 461535 4029
rect 509249 3995 509283 4777
rect 509341 4131 509375 4777
rect 504465 3655 504499 3961
rect 513941 3655 513975 4097
rect 514033 3927 514067 4097
rect 514125 3723 514159 3893
rect 516149 3723 516183 3961
rect 514217 3655 514251 3689
rect 513941 3621 514251 3655
rect 521945 3519 521979 5525
rect 523601 3519 523635 3553
rect 523601 3485 523785 3519
rect 461075 3009 461351 3043
rect 518909 2635 518943 3417
<< viali >>
rect 292497 11033 292531 11067
rect 282837 10965 282871 10999
rect 292313 10965 292347 10999
rect 292405 10965 292439 10999
rect 302249 10965 302283 10999
rect 277593 10761 277627 10795
rect 286885 10761 286919 10795
rect 287253 10557 287287 10591
rect 287621 10557 287655 10591
rect 302249 10761 302283 10795
rect 287805 10489 287839 10523
rect 292313 10489 292347 10523
rect 278145 10421 278179 10455
rect 282745 10421 282779 10455
rect 307217 10693 307251 10727
rect 306389 10557 306423 10591
rect 302433 10489 302467 10523
rect 306205 10489 306239 10523
rect 306941 10557 306975 10591
rect 302249 10149 302283 10183
rect 302341 10149 302375 10183
rect 311633 10625 311667 10659
rect 311541 10557 311575 10591
rect 311909 10557 311943 10591
rect 311817 10489 311851 10523
rect 307217 10149 307251 10183
rect 307309 10149 307343 10183
rect 307125 10013 307159 10047
rect 306941 9945 306975 9979
rect 302249 9605 302283 9639
rect 284125 9469 284159 9503
rect 292497 9469 292531 9503
rect 284401 9333 284435 9367
rect 287529 9333 287563 9367
rect 287621 9333 287655 9367
rect 292313 9129 292347 9163
rect 292497 9129 292531 9163
rect 287621 9061 287655 9095
rect 287805 8993 287839 9027
rect 292405 8993 292439 9027
rect 292497 8993 292531 9027
rect 253213 8245 253247 8279
rect 253213 8041 253247 8075
rect 253305 8041 253339 8075
rect 253305 7701 253339 7735
rect 253489 7769 253523 7803
rect 253489 7361 253523 7395
rect 292497 7361 292531 7395
rect 463893 7497 463927 7531
rect 400045 7293 400079 7327
rect 400321 7157 400355 7191
rect 398113 6749 398147 6783
rect 348893 6681 348927 6715
rect 394525 6613 394559 6647
rect 398021 6613 398055 6647
rect 398113 6613 398147 6647
rect 398205 6749 398239 6783
rect 349353 6409 349387 6443
rect 394433 6409 394467 6443
rect 394525 6409 394559 6443
rect 349905 6273 349939 6307
rect 394801 6273 394835 6307
rect 327733 5797 327767 5831
rect 320741 5661 320775 5695
rect 209421 5593 209455 5627
rect 219633 5593 219667 5627
rect 209421 5253 209455 5287
rect 209513 5525 209547 5559
rect 209513 5185 209547 5219
rect 209605 5253 209639 5287
rect 209697 5185 209731 5219
rect 277041 5593 277075 5627
rect 219725 5525 219759 5559
rect 465825 7497 465859 7531
rect 465733 7361 465767 7395
rect 465733 6885 465767 6919
rect 465825 6885 465859 6919
rect 502257 6885 502291 6919
rect 349905 5593 349939 5627
rect 388453 6205 388487 6239
rect 277041 5321 277075 5355
rect 279709 5525 279743 5559
rect 278237 5253 278271 5287
rect 278421 5253 278455 5287
rect 282653 5525 282687 5559
rect 320649 5525 320683 5559
rect 320741 5525 320775 5559
rect 321017 5525 321051 5559
rect 327733 5525 327767 5559
rect 463709 6205 463743 6239
rect 463893 6205 463927 6239
rect 463985 6205 464019 6239
rect 502257 6137 502291 6171
rect 388453 5525 388487 5559
rect 509341 5525 509375 5559
rect 282653 5321 282687 5355
rect 219725 5117 219759 5151
rect 278145 5185 278179 5219
rect 279709 5185 279743 5219
rect 209513 4981 209547 5015
rect 219541 5049 219575 5083
rect 219633 5049 219667 5083
rect 209421 4777 209455 4811
rect 123217 4165 123251 4199
rect 116317 3689 116351 3723
rect 34529 3553 34563 3587
rect 34529 3349 34563 3383
rect 92489 3349 92523 3383
rect 92489 3145 92523 3179
rect 116317 2805 116351 2839
rect 128553 4165 128587 4199
rect 124597 3689 124631 3723
rect 127633 3621 127667 3655
rect 124597 3485 124631 3519
rect 126897 3485 126931 3519
rect 123217 2805 123251 2839
rect 123309 3417 123343 3451
rect 123309 2805 123343 2839
rect 127541 3417 127575 3451
rect 127633 3417 127667 3451
rect 127725 3621 127759 3655
rect 128553 3621 128587 3655
rect 132785 4165 132819 4199
rect 277869 4709 277903 4743
rect 278053 4641 278087 4675
rect 509341 4981 509375 5015
rect 521945 5525 521979 5559
rect 278145 4573 278179 4607
rect 509249 4777 509283 4811
rect 219541 4097 219575 4131
rect 461317 4097 461351 4131
rect 128461 3485 128495 3519
rect 132785 3485 132819 3519
rect 132877 4029 132911 4063
rect 461041 4029 461075 4063
rect 451289 3893 451323 3927
rect 451381 3689 451415 3723
rect 455429 3893 455463 3927
rect 455429 3689 455463 3723
rect 460765 3893 460799 3927
rect 426081 3621 426115 3655
rect 132877 3485 132911 3519
rect 156981 3485 157015 3519
rect 128645 3417 128679 3451
rect 158545 3417 158579 3451
rect 158729 3417 158763 3451
rect 156981 3349 157015 3383
rect 426081 2941 426115 2975
rect 126897 2601 126931 2635
rect 128461 2805 128495 2839
rect 132325 2805 132359 2839
rect 436661 2805 436695 2839
rect 437489 2805 437523 2839
rect 132325 2601 132359 2635
rect 460949 3349 460983 3383
rect 461041 3349 461075 3383
rect 461225 3077 461259 3111
rect 462513 4029 462547 4063
rect 509341 4777 509375 4811
rect 509341 4097 509375 4131
rect 513941 4097 513975 4131
rect 504465 3961 504499 3995
rect 509249 3961 509283 3995
rect 504465 3621 504499 3655
rect 514033 4097 514067 4131
rect 516149 3961 516183 3995
rect 514033 3893 514067 3927
rect 514125 3893 514159 3927
rect 514125 3689 514159 3723
rect 514217 3689 514251 3723
rect 516149 3689 516183 3723
rect 521945 3485 521979 3519
rect 523601 3553 523635 3587
rect 523785 3485 523819 3519
rect 461501 3417 461535 3451
rect 518909 3417 518943 3451
rect 461041 3009 461075 3043
rect 460765 2601 460799 2635
rect 518909 2601 518943 2635
rect 128461 2533 128495 2567
<< metal1 >>
rect 1104 701712 582820 701808
rect 1104 701168 582820 701264
rect 1104 700624 582820 700720
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 41322 700516 41328 700528
rect 40552 700488 41328 700516
rect 40552 700476 40558 700488
rect 41322 700476 41328 700488
rect 41380 700476 41386 700528
rect 480162 700476 480168 700528
rect 480220 700516 480226 700528
rect 527174 700516 527180 700528
rect 480220 700488 527180 700516
rect 480220 700476 480226 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 402882 700408 402888 700460
rect 402940 700448 402946 700460
rect 429838 700448 429844 700460
rect 402940 700420 429844 700448
rect 402940 700408 402946 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 441522 700408 441528 700460
rect 441580 700448 441586 700460
rect 478506 700448 478512 700460
rect 441580 700420 478512 700448
rect 441580 700408 441586 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 492582 700408 492588 700460
rect 492640 700448 492646 700460
rect 543458 700448 543464 700460
rect 492640 700420 543464 700448
rect 492640 700408 492646 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 378042 700340 378048 700392
rect 378100 700380 378106 700392
rect 397454 700380 397460 700392
rect 378100 700352 397460 700380
rect 378100 700340 378106 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 416682 700340 416688 700392
rect 416740 700380 416746 700392
rect 446122 700380 446128 700392
rect 416740 700352 446128 700380
rect 416740 700340 416746 700352
rect 446122 700340 446128 700352
rect 446180 700340 446186 700392
rect 453942 700340 453948 700392
rect 454000 700380 454006 700392
rect 494790 700380 494796 700392
rect 454000 700352 494796 700380
rect 454000 700340 454006 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 506382 700340 506388 700392
rect 506440 700380 506446 700392
rect 559650 700380 559656 700392
rect 506440 700352 559656 700380
rect 506440 700340 506446 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 56778 700272 56784 700324
rect 56836 700312 56842 700324
rect 57882 700312 57888 700324
rect 56836 700284 57888 700312
rect 56836 700272 56842 700284
rect 57882 700272 57888 700284
rect 57940 700272 57946 700324
rect 186498 700272 186504 700324
rect 186556 700312 186562 700324
rect 187602 700312 187608 700324
rect 186556 700284 187608 700312
rect 186556 700272 186562 700284
rect 187602 700272 187608 700284
rect 187660 700272 187666 700324
rect 339402 700272 339408 700324
rect 339460 700312 339466 700324
rect 348786 700312 348792 700324
rect 339460 700284 348792 700312
rect 339460 700272 339466 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 351822 700272 351828 700324
rect 351880 700312 351886 700324
rect 364978 700312 364984 700324
rect 351880 700284 364984 700312
rect 351880 700272 351886 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 365622 700272 365628 700324
rect 365680 700312 365686 700324
rect 381170 700312 381176 700324
rect 365680 700284 381176 700312
rect 365680 700272 365686 700284
rect 381170 700272 381176 700284
rect 381228 700272 381234 700324
rect 390462 700272 390468 700324
rect 390520 700312 390526 700324
rect 413646 700312 413652 700324
rect 390520 700284 413652 700312
rect 390520 700272 390526 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 467742 700272 467748 700324
rect 467800 700312 467806 700324
rect 510982 700312 510988 700324
rect 467800 700284 510988 700312
rect 467800 700272 467806 700284
rect 510982 700272 510988 700284
rect 511040 700272 511046 700324
rect 517422 700272 517428 700324
rect 517480 700312 517486 700324
rect 575842 700312 575848 700324
rect 517480 700284 575848 700312
rect 517480 700272 517486 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 1104 700080 582820 700176
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 251450 699660 251456 699712
rect 251508 699700 251514 699712
rect 252462 699700 252468 699712
rect 251508 699672 252468 699700
rect 251508 699660 251514 699672
rect 252462 699660 252468 699672
rect 252520 699660 252526 699712
rect 299474 699660 299480 699712
rect 299532 699700 299538 699712
rect 300118 699700 300124 699712
rect 299532 699672 300124 699700
rect 299532 699660 299538 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 313182 699660 313188 699712
rect 313240 699700 313246 699712
rect 316310 699700 316316 699712
rect 313240 699672 316316 699700
rect 313240 699660 313246 699672
rect 316310 699660 316316 699672
rect 316368 699660 316374 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 332502 699700 332508 699712
rect 327040 699672 332508 699700
rect 327040 699660 327046 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 1104 699536 582820 699632
rect 1104 698992 582820 699088
rect 1104 698448 582820 698544
rect 1104 697904 582820 698000
rect 1104 697360 582820 697456
rect 520918 696940 520924 696992
rect 520976 696980 520982 696992
rect 580166 696980 580172 696992
rect 520976 696952 580172 696980
rect 520976 696940 520982 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 1104 696816 582820 696912
rect 1104 696272 582820 696368
rect 1104 695728 582820 695824
rect 1104 695184 582820 695280
rect 1104 694640 582820 694736
rect 1104 694096 582820 694192
rect 1104 693552 582820 693648
rect 1104 693008 582820 693104
rect 1104 692464 582820 692560
rect 1104 691920 582820 692016
rect 1104 691376 582820 691472
rect 1104 690832 582820 690928
rect 1104 690288 582820 690384
rect 1104 689744 582820 689840
rect 1104 689200 582820 689296
rect 1104 688656 582820 688752
rect 1104 688112 582820 688208
rect 1104 687568 582820 687664
rect 1104 687024 582820 687120
rect 1104 686480 582820 686576
rect 1104 685936 582820 686032
rect 1104 685392 582820 685488
rect 1104 684848 582820 684944
rect 1104 684304 582820 684400
rect 1104 683760 582820 683856
rect 1104 683216 582820 683312
rect 521010 683136 521016 683188
rect 521068 683176 521074 683188
rect 580166 683176 580172 683188
rect 521068 683148 580172 683176
rect 521068 683136 521074 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 284202 682864 284208 682916
rect 284260 682904 284266 682916
rect 287606 682904 287612 682916
rect 284260 682876 287612 682904
rect 284260 682864 284266 682876
rect 287606 682864 287612 682876
rect 287664 682864 287670 682916
rect 1104 682672 582820 682768
rect 57882 682592 57888 682644
rect 57940 682632 57946 682644
rect 108390 682632 108396 682644
rect 57940 682604 108396 682632
rect 57940 682592 57946 682604
rect 108390 682592 108396 682604
rect 108448 682592 108454 682644
rect 41322 682524 41328 682576
rect 41380 682564 41386 682576
rect 95602 682564 95608 682576
rect 41380 682536 95608 682564
rect 41380 682524 41386 682536
rect 95602 682524 95608 682536
rect 95660 682524 95666 682576
rect 106182 682524 106188 682576
rect 106240 682564 106246 682576
rect 146846 682564 146852 682576
rect 106240 682536 146852 682564
rect 106240 682524 106246 682536
rect 146846 682524 146852 682536
rect 146904 682524 146910 682576
rect 154482 682524 154488 682576
rect 154540 682564 154546 682576
rect 185210 682564 185216 682576
rect 154540 682536 185216 682564
rect 154540 682524 154546 682536
rect 185210 682524 185216 682536
rect 185268 682524 185274 682576
rect 24762 682456 24768 682508
rect 24820 682496 24826 682508
rect 82814 682496 82820 682508
rect 24820 682468 82820 682496
rect 24820 682456 24826 682468
rect 82814 682456 82820 682468
rect 82872 682456 82878 682508
rect 89622 682456 89628 682508
rect 89680 682496 89686 682508
rect 134058 682496 134064 682508
rect 89680 682468 134064 682496
rect 89680 682456 89686 682468
rect 134058 682456 134064 682468
rect 134116 682456 134122 682508
rect 137922 682456 137928 682508
rect 137980 682496 137986 682508
rect 172422 682496 172428 682508
rect 137980 682468 172428 682496
rect 137980 682456 137986 682468
rect 172422 682456 172428 682468
rect 172480 682456 172486 682508
rect 187602 682456 187608 682508
rect 187660 682496 187666 682508
rect 210786 682496 210792 682508
rect 187660 682468 210792 682496
rect 187660 682456 187666 682468
rect 210786 682456 210792 682468
rect 210844 682456 210850 682508
rect 219342 682456 219348 682508
rect 219400 682496 219406 682508
rect 236362 682496 236368 682508
rect 219400 682468 236368 682496
rect 219400 682456 219406 682468
rect 236362 682456 236368 682468
rect 236420 682456 236426 682508
rect 8202 682388 8208 682440
rect 8260 682428 8266 682440
rect 71038 682428 71044 682440
rect 8260 682400 71044 682428
rect 8260 682388 8266 682400
rect 71038 682388 71044 682400
rect 71096 682388 71102 682440
rect 73062 682388 73068 682440
rect 73120 682428 73126 682440
rect 121178 682428 121184 682440
rect 73120 682400 121184 682428
rect 73120 682388 73126 682400
rect 121178 682388 121184 682400
rect 121236 682388 121242 682440
rect 122742 682388 122748 682440
rect 122800 682428 122806 682440
rect 159634 682428 159640 682440
rect 122800 682400 159640 682428
rect 122800 682388 122806 682400
rect 159634 682388 159640 682400
rect 159692 682388 159698 682440
rect 171042 682388 171048 682440
rect 171100 682428 171106 682440
rect 197998 682428 198004 682440
rect 171100 682400 198004 682428
rect 171100 682388 171106 682400
rect 197998 682388 198004 682400
rect 198056 682388 198062 682440
rect 202782 682388 202788 682440
rect 202840 682428 202846 682440
rect 223574 682428 223580 682440
rect 202840 682400 223580 682428
rect 202840 682388 202846 682400
rect 223574 682388 223580 682400
rect 223632 682388 223638 682440
rect 235902 682388 235908 682440
rect 235960 682428 235966 682440
rect 249242 682428 249248 682440
rect 235960 682400 249248 682428
rect 235960 682388 235966 682400
rect 249242 682388 249248 682400
rect 249300 682388 249306 682440
rect 252462 682388 252468 682440
rect 252520 682428 252526 682440
rect 262030 682428 262036 682440
rect 252520 682400 262036 682428
rect 252520 682388 252526 682400
rect 262030 682388 262036 682400
rect 262088 682388 262094 682440
rect 267642 682388 267648 682440
rect 267700 682428 267706 682440
rect 274818 682428 274824 682440
rect 267700 682400 274824 682428
rect 267700 682388 267706 682400
rect 274818 682388 274824 682400
rect 274876 682388 274882 682440
rect 1104 682128 582820 682224
rect 325970 681708 325976 681760
rect 326028 681748 326034 681760
rect 326982 681748 326988 681760
rect 326028 681720 326988 681748
rect 326028 681708 326034 681720
rect 326982 681708 326988 681720
rect 327040 681708 327046 681760
rect 338758 681708 338764 681760
rect 338816 681748 338822 681760
rect 339402 681748 339408 681760
rect 338816 681720 339408 681748
rect 338816 681708 338822 681720
rect 339402 681708 339408 681720
rect 339460 681708 339466 681760
rect 364426 681708 364432 681760
rect 364484 681748 364490 681760
rect 365622 681748 365628 681760
rect 364484 681720 365628 681748
rect 364484 681708 364490 681720
rect 365622 681708 365628 681720
rect 365680 681708 365686 681760
rect 377214 681708 377220 681760
rect 377272 681748 377278 681760
rect 378042 681748 378048 681760
rect 377272 681720 378048 681748
rect 377272 681708 377278 681720
rect 378042 681708 378048 681720
rect 378100 681708 378106 681760
rect 390002 681708 390008 681760
rect 390060 681748 390066 681760
rect 390462 681748 390468 681760
rect 390060 681720 390468 681748
rect 390060 681708 390066 681720
rect 390462 681708 390468 681720
rect 390520 681708 390526 681760
rect 415578 681708 415584 681760
rect 415636 681748 415642 681760
rect 416682 681748 416688 681760
rect 415636 681720 416688 681748
rect 415636 681708 415642 681720
rect 416682 681708 416688 681720
rect 416740 681708 416746 681760
rect 428366 681708 428372 681760
rect 428424 681748 428430 681760
rect 429102 681748 429108 681760
rect 428424 681720 429108 681748
rect 428424 681708 428430 681720
rect 429102 681708 429108 681720
rect 429160 681708 429166 681760
rect 466730 681708 466736 681760
rect 466788 681748 466794 681760
rect 467742 681748 467748 681760
rect 466788 681720 467748 681748
rect 466788 681708 466794 681720
rect 467742 681708 467748 681720
rect 467800 681708 467806 681760
rect 479610 681708 479616 681760
rect 479668 681748 479674 681760
rect 480162 681748 480168 681760
rect 479668 681720 480168 681748
rect 479668 681708 479674 681720
rect 480162 681708 480168 681720
rect 480220 681708 480226 681760
rect 505186 681708 505192 681760
rect 505244 681748 505250 681760
rect 506382 681748 506388 681760
rect 505244 681720 506388 681748
rect 505244 681708 505250 681720
rect 506382 681708 506388 681720
rect 506440 681708 506446 681760
rect 1104 681584 68000 681680
rect 519948 681584 582820 681680
rect 1104 681040 68000 681136
rect 519948 681040 582820 681136
rect 1104 680496 68000 680592
rect 519948 680496 582820 680592
rect 3418 680280 3424 680332
rect 3476 680320 3482 680332
rect 66990 680320 66996 680332
rect 3476 680292 66996 680320
rect 3476 680280 3482 680292
rect 66990 680280 66996 680292
rect 67048 680280 67054 680332
rect 1104 679952 68000 680048
rect 519948 679952 582820 680048
rect 1104 679408 68000 679504
rect 519948 679408 582820 679504
rect 1104 678864 68000 678960
rect 519948 678864 582820 678960
rect 1104 678320 68000 678416
rect 519948 678320 582820 678416
rect 1104 677776 68000 677872
rect 519948 677776 582820 677872
rect 1104 677232 68000 677328
rect 519948 677232 582820 677328
rect 1104 676688 68000 676784
rect 519948 676688 582820 676784
rect 1104 676144 68000 676240
rect 519948 676144 582820 676240
rect 1104 675600 68000 675696
rect 519948 675600 582820 675696
rect 1104 675056 68000 675152
rect 519948 675056 582820 675152
rect 1104 674512 68000 674608
rect 519948 674512 582820 674608
rect 1104 673968 68000 674064
rect 519948 673968 582820 674064
rect 1104 673424 68000 673520
rect 519948 673424 582820 673520
rect 1104 672880 68000 672976
rect 519948 672880 582820 672976
rect 1104 672336 68000 672432
rect 519948 672336 582820 672432
rect 1104 671792 68000 671888
rect 519948 671792 582820 671888
rect 1104 671248 68000 671344
rect 519948 671248 582820 671344
rect 520918 670828 520924 670880
rect 520976 670868 520982 670880
rect 580166 670868 580172 670880
rect 520976 670840 580172 670868
rect 520976 670828 520982 670840
rect 580166 670828 580172 670840
rect 580224 670828 580230 670880
rect 1104 670704 68000 670800
rect 519948 670704 582820 670800
rect 1104 670160 68000 670256
rect 519948 670160 582820 670256
rect 1104 669616 68000 669712
rect 519948 669616 582820 669712
rect 3510 669264 3516 669316
rect 3568 669304 3574 669316
rect 67174 669304 67180 669316
rect 3568 669276 67180 669304
rect 3568 669264 3574 669276
rect 67174 669264 67180 669276
rect 67232 669264 67238 669316
rect 1104 669072 68000 669168
rect 519948 669072 582820 669168
rect 1104 668528 68000 668624
rect 519948 668528 582820 668624
rect 1104 667984 68000 668080
rect 519948 667984 582820 668080
rect 1104 667440 68000 667536
rect 519948 667440 582820 667536
rect 1104 666896 68000 666992
rect 519948 666896 582820 666992
rect 1104 666352 68000 666448
rect 519948 666352 582820 666448
rect 1104 665808 68000 665904
rect 519948 665808 582820 665904
rect 1104 665264 68000 665360
rect 519948 665264 582820 665360
rect 1104 664720 68000 664816
rect 519948 664720 582820 664816
rect 1104 664176 68000 664272
rect 519948 664176 582820 664272
rect 1104 663632 68000 663728
rect 519948 663632 582820 663728
rect 1104 663088 68000 663184
rect 519948 663088 582820 663184
rect 1104 662544 68000 662640
rect 519948 662544 582820 662640
rect 1104 662000 68000 662096
rect 519948 662000 582820 662096
rect 1104 661456 68000 661552
rect 519948 661456 582820 661552
rect 1104 660912 68000 661008
rect 519948 660912 582820 661008
rect 1104 660368 68000 660464
rect 519948 660368 582820 660464
rect 1104 659824 68000 659920
rect 519948 659824 582820 659920
rect 1104 659280 68000 659376
rect 519948 659280 582820 659376
rect 1104 658736 68000 658832
rect 519948 658736 582820 658832
rect 1104 658192 68000 658288
rect 519948 658192 582820 658288
rect 3418 658112 3424 658164
rect 3476 658152 3482 658164
rect 67358 658152 67364 658164
rect 3476 658124 67364 658152
rect 3476 658112 3482 658124
rect 67358 658112 67364 658124
rect 67416 658112 67422 658164
rect 1104 657648 68000 657744
rect 519948 657648 582820 657744
rect 1104 657104 68000 657200
rect 519948 657104 582820 657200
rect 521010 656888 521016 656940
rect 521068 656928 521074 656940
rect 580166 656928 580172 656940
rect 521068 656900 580172 656928
rect 521068 656888 521074 656900
rect 580166 656888 580172 656900
rect 580224 656888 580230 656940
rect 1104 656560 68000 656656
rect 519948 656560 582820 656656
rect 1104 656016 68000 656112
rect 519948 656016 582820 656112
rect 1104 655472 68000 655568
rect 519948 655472 582820 655568
rect 1104 654928 68000 655024
rect 519948 654928 582820 655024
rect 1104 654384 68000 654480
rect 519948 654384 582820 654480
rect 1104 653840 68000 653936
rect 519948 653840 582820 653936
rect 1104 653296 68000 653392
rect 519948 653296 582820 653392
rect 1104 652752 68000 652848
rect 519948 652752 582820 652848
rect 1104 652208 68000 652304
rect 519948 652208 582820 652304
rect 1104 651664 68000 651760
rect 519948 651664 582820 651760
rect 1104 651120 68000 651216
rect 519948 651120 582820 651216
rect 1104 650576 68000 650672
rect 519948 650576 582820 650672
rect 1104 650032 68000 650128
rect 519948 650032 582820 650128
rect 1104 649488 68000 649584
rect 519948 649488 582820 649584
rect 1104 648944 68000 649040
rect 519948 648944 582820 649040
rect 1104 648400 68000 648496
rect 519948 648400 582820 648496
rect 1104 647856 68000 647952
rect 519948 647856 582820 647952
rect 1104 647312 68000 647408
rect 519948 647312 582820 647408
rect 3510 647164 3516 647216
rect 3568 647204 3574 647216
rect 67358 647204 67364 647216
rect 3568 647176 67364 647204
rect 3568 647164 3574 647176
rect 67358 647164 67364 647176
rect 67416 647164 67422 647216
rect 1104 646768 68000 646864
rect 519948 646768 582820 646864
rect 1104 646224 68000 646320
rect 519948 646224 582820 646320
rect 1104 645680 68000 645776
rect 519948 645680 582820 645776
rect 1104 645136 68000 645232
rect 519948 645136 582820 645232
rect 1104 644592 68000 644688
rect 519948 644592 582820 644688
rect 1104 644048 68000 644144
rect 519948 644048 582820 644144
rect 1104 643504 68000 643600
rect 519948 643504 582820 643600
rect 520918 643084 520924 643136
rect 520976 643124 520982 643136
rect 580166 643124 580172 643136
rect 520976 643096 580172 643124
rect 520976 643084 520982 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 1104 642960 68000 643056
rect 519948 642960 582820 643056
rect 1104 642416 68000 642512
rect 519948 642416 582820 642512
rect 1104 641872 68000 641968
rect 519948 641872 582820 641968
rect 1104 641328 68000 641424
rect 519948 641328 582820 641424
rect 1104 640784 68000 640880
rect 519948 640784 582820 640880
rect 1104 640240 68000 640336
rect 519948 640240 582820 640336
rect 1104 639696 68000 639792
rect 519948 639696 582820 639792
rect 1104 639152 68000 639248
rect 519948 639152 582820 639248
rect 1104 638608 68000 638704
rect 519948 638608 582820 638704
rect 1104 638064 68000 638160
rect 519948 638064 582820 638160
rect 1104 637520 68000 637616
rect 519948 637520 582820 637616
rect 1104 636976 68000 637072
rect 519948 636976 582820 637072
rect 1104 636432 68000 636528
rect 519948 636432 582820 636528
rect 3418 636148 3424 636200
rect 3476 636188 3482 636200
rect 67358 636188 67364 636200
rect 3476 636160 67364 636188
rect 3476 636148 3482 636160
rect 67358 636148 67364 636160
rect 67416 636148 67422 636200
rect 1104 635888 68000 635984
rect 519948 635888 582820 635984
rect 1104 635344 68000 635440
rect 519948 635344 582820 635440
rect 1104 634800 68000 634896
rect 519948 634800 582820 634896
rect 1104 634256 68000 634352
rect 519948 634256 582820 634352
rect 1104 633712 68000 633808
rect 519948 633712 582820 633808
rect 1104 633168 68000 633264
rect 519948 633168 582820 633264
rect 1104 632624 68000 632720
rect 519948 632624 582820 632720
rect 1104 632080 68000 632176
rect 519948 632080 582820 632176
rect 1104 631536 68000 631632
rect 519948 631536 582820 631632
rect 1104 630992 68000 631088
rect 519948 630992 582820 631088
rect 520918 630640 520924 630692
rect 520976 630680 520982 630692
rect 580166 630680 580172 630692
rect 520976 630652 580172 630680
rect 520976 630640 520982 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 1104 630448 68000 630544
rect 519948 630448 582820 630544
rect 1104 629904 68000 630000
rect 519948 629904 582820 630000
rect 1104 629360 68000 629456
rect 519948 629360 582820 629456
rect 1104 628816 68000 628912
rect 519948 628816 582820 628912
rect 1104 628272 68000 628368
rect 519948 628272 582820 628368
rect 1104 627728 68000 627824
rect 519948 627728 582820 627824
rect 1104 627184 68000 627280
rect 519948 627184 582820 627280
rect 1104 626640 68000 626736
rect 519948 626640 582820 626736
rect 1104 626096 68000 626192
rect 519948 626096 582820 626192
rect 1104 625552 68000 625648
rect 519948 625552 582820 625648
rect 1104 625008 68000 625104
rect 519948 625008 582820 625104
rect 3418 624928 3424 624980
rect 3476 624968 3482 624980
rect 67358 624968 67364 624980
rect 3476 624940 67364 624968
rect 3476 624928 3482 624940
rect 67358 624928 67364 624940
rect 67416 624928 67422 624980
rect 1104 624464 68000 624560
rect 519948 624464 582820 624560
rect 1104 623920 68000 624016
rect 519948 623920 582820 624016
rect 1104 623376 68000 623472
rect 519948 623376 582820 623472
rect 1104 622832 68000 622928
rect 519948 622832 582820 622928
rect 1104 622288 68000 622384
rect 519948 622288 582820 622384
rect 1104 621744 68000 621840
rect 519948 621744 582820 621840
rect 1104 621200 68000 621296
rect 519948 621200 582820 621296
rect 1104 620656 68000 620752
rect 519948 620656 582820 620752
rect 1104 620112 68000 620208
rect 519948 620112 582820 620208
rect 1104 619568 68000 619664
rect 519948 619568 582820 619664
rect 1104 619024 68000 619120
rect 519948 619024 582820 619120
rect 1104 618480 68000 618576
rect 519948 618480 582820 618576
rect 1104 617936 68000 618032
rect 519948 617936 582820 618032
rect 1104 617392 68000 617488
rect 519948 617392 582820 617488
rect 520274 616972 520280 617024
rect 520332 617012 520338 617024
rect 580166 617012 580172 617024
rect 520332 616984 580172 617012
rect 520332 616972 520338 616984
rect 580166 616972 580172 616984
rect 580224 616972 580230 617024
rect 1104 616848 68000 616944
rect 519948 616848 582820 616944
rect 1104 616304 68000 616400
rect 519948 616304 582820 616400
rect 1104 615760 68000 615856
rect 519948 615760 582820 615856
rect 1104 615216 68000 615312
rect 519948 615216 582820 615312
rect 1104 614672 68000 614768
rect 519948 614672 582820 614768
rect 1104 614128 68000 614224
rect 519948 614128 582820 614224
rect 3418 614048 3424 614100
rect 3476 614088 3482 614100
rect 66898 614088 66904 614100
rect 3476 614060 66904 614088
rect 3476 614048 3482 614060
rect 66898 614048 66904 614060
rect 66956 614048 66962 614100
rect 1104 613584 68000 613680
rect 519948 613584 582820 613680
rect 1104 613040 68000 613136
rect 519948 613040 582820 613136
rect 1104 612496 68000 612592
rect 519948 612496 582820 612592
rect 1104 611952 68000 612048
rect 519948 611952 582820 612048
rect 1104 611408 68000 611504
rect 519948 611408 582820 611504
rect 1104 610864 68000 610960
rect 519948 610864 582820 610960
rect 1104 610320 68000 610416
rect 519948 610320 582820 610416
rect 1104 609776 68000 609872
rect 519948 609776 582820 609872
rect 1104 609232 68000 609328
rect 519948 609232 582820 609328
rect 1104 608688 68000 608784
rect 519948 608688 582820 608784
rect 1104 608144 68000 608240
rect 519948 608144 582820 608240
rect 1104 607600 68000 607696
rect 519948 607600 582820 607696
rect 1104 607056 68000 607152
rect 519948 607056 582820 607152
rect 1104 606512 68000 606608
rect 519948 606512 582820 606608
rect 1104 605968 68000 606064
rect 519948 605968 582820 606064
rect 1104 605424 68000 605520
rect 519948 605424 582820 605520
rect 1104 604880 68000 604976
rect 519948 604880 582820 604976
rect 1104 604336 68000 604432
rect 519948 604336 582820 604432
rect 1104 603792 68000 603888
rect 519948 603792 582820 603888
rect 1104 603248 68000 603344
rect 519948 603248 582820 603344
rect 521102 603100 521108 603152
rect 521160 603140 521166 603152
rect 580166 603140 580172 603152
rect 521160 603112 580172 603140
rect 521160 603100 521166 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 4062 603032 4068 603084
rect 4120 603072 4126 603084
rect 66438 603072 66444 603084
rect 4120 603044 66444 603072
rect 4120 603032 4126 603044
rect 66438 603032 66444 603044
rect 66496 603032 66502 603084
rect 1104 602704 68000 602800
rect 519948 602704 582820 602800
rect 1104 602160 68000 602256
rect 519948 602160 582820 602256
rect 1104 601616 68000 601712
rect 519948 601616 582820 601712
rect 1104 601072 68000 601168
rect 519948 601072 582820 601168
rect 1104 600528 68000 600624
rect 519948 600528 582820 600624
rect 1104 599984 68000 600080
rect 519948 599984 582820 600080
rect 1104 599440 68000 599536
rect 519948 599440 582820 599536
rect 1104 598896 68000 598992
rect 519948 598896 582820 598992
rect 1104 598352 68000 598448
rect 519948 598352 582820 598448
rect 1104 597808 68000 597904
rect 519948 597808 582820 597904
rect 1104 597264 68000 597360
rect 519948 597264 582820 597360
rect 1104 596720 68000 596816
rect 519948 596720 582820 596816
rect 1104 596176 68000 596272
rect 519948 596176 582820 596272
rect 1104 595632 68000 595728
rect 519948 595632 582820 595728
rect 1104 595088 68000 595184
rect 519948 595088 582820 595184
rect 1104 594544 68000 594640
rect 519948 594544 582820 594640
rect 1104 594000 68000 594096
rect 519948 594000 582820 594096
rect 1104 593456 68000 593552
rect 519948 593456 582820 593552
rect 1104 592912 68000 593008
rect 519948 592912 582820 593008
rect 1104 592368 68000 592464
rect 519948 592368 582820 592464
rect 3418 591948 3424 592000
rect 3476 591988 3482 592000
rect 66990 591988 66996 592000
rect 3476 591960 66996 591988
rect 3476 591948 3482 591960
rect 66990 591948 66996 591960
rect 67048 591948 67054 592000
rect 1104 591824 68000 591920
rect 519948 591824 582820 591920
rect 1104 591280 68000 591376
rect 519948 591280 582820 591376
rect 1104 590736 68000 590832
rect 519948 590736 582820 590832
rect 521562 590656 521568 590708
rect 521620 590696 521626 590708
rect 579798 590696 579804 590708
rect 521620 590668 579804 590696
rect 521620 590656 521626 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 1104 590192 68000 590288
rect 519948 590192 582820 590288
rect 1104 589648 68000 589744
rect 519948 589648 582820 589744
rect 1104 589104 68000 589200
rect 519948 589104 582820 589200
rect 1104 588560 68000 588656
rect 519948 588560 582820 588656
rect 1104 588016 68000 588112
rect 519948 588016 582820 588112
rect 1104 587472 68000 587568
rect 519948 587472 582820 587568
rect 1104 586928 68000 587024
rect 519948 586928 582820 587024
rect 1104 586384 68000 586480
rect 519948 586384 582820 586480
rect 1104 585840 68000 585936
rect 519948 585840 582820 585936
rect 1104 585296 68000 585392
rect 519948 585296 582820 585392
rect 1104 584752 68000 584848
rect 519948 584752 582820 584848
rect 1104 584208 68000 584304
rect 519948 584208 582820 584304
rect 1104 583664 68000 583760
rect 519948 583664 582820 583760
rect 1104 583120 68000 583216
rect 519948 583120 582820 583216
rect 1104 582576 68000 582672
rect 519948 582576 582820 582672
rect 1104 582032 68000 582128
rect 519948 582032 582820 582128
rect 1104 581488 68000 581584
rect 519948 581488 582820 581584
rect 1104 580944 68000 581040
rect 519948 580944 582820 581040
rect 1104 580400 68000 580496
rect 519948 580400 582820 580496
rect 1104 579856 68000 579952
rect 519948 579856 582820 579952
rect 3418 579572 3424 579624
rect 3476 579612 3482 579624
rect 67174 579612 67180 579624
rect 3476 579584 67180 579612
rect 3476 579572 3482 579584
rect 67174 579572 67180 579584
rect 67232 579572 67238 579624
rect 1104 579312 68000 579408
rect 519948 579312 582820 579408
rect 1104 578768 68000 578864
rect 519948 578768 582820 578864
rect 1104 578224 68000 578320
rect 519948 578224 582820 578320
rect 1104 577680 68000 577776
rect 519948 577680 582820 577776
rect 521562 577464 521568 577516
rect 521620 577504 521626 577516
rect 580166 577504 580172 577516
rect 521620 577476 580172 577504
rect 521620 577464 521626 577476
rect 580166 577464 580172 577476
rect 580224 577464 580230 577516
rect 1104 577136 68000 577232
rect 519948 577136 582820 577232
rect 1104 576592 68000 576688
rect 519948 576592 582820 576688
rect 1104 576048 68000 576144
rect 519948 576048 582820 576144
rect 1104 575504 68000 575600
rect 519948 575504 582820 575600
rect 1104 574960 68000 575056
rect 519948 574960 582820 575056
rect 1104 574416 68000 574512
rect 519948 574416 582820 574512
rect 1104 573872 68000 573968
rect 519948 573872 582820 573968
rect 1104 573328 68000 573424
rect 519948 573328 582820 573424
rect 1104 572784 68000 572880
rect 519948 572784 582820 572880
rect 1104 572240 68000 572336
rect 519948 572240 582820 572336
rect 1104 571696 68000 571792
rect 519948 571696 582820 571792
rect 1104 571152 68000 571248
rect 519948 571152 582820 571248
rect 1104 570608 68000 570704
rect 519948 570608 582820 570704
rect 1104 570064 68000 570160
rect 519948 570064 582820 570160
rect 1104 569520 68000 569616
rect 519948 569520 582820 569616
rect 1104 568976 68000 569072
rect 519948 568976 582820 569072
rect 1104 568432 68000 568528
rect 519948 568432 582820 568528
rect 1104 567888 68000 567984
rect 519948 567888 582820 567984
rect 1104 567344 68000 567440
rect 519948 567344 582820 567440
rect 4062 567196 4068 567248
rect 4120 567236 4126 567248
rect 67358 567236 67364 567248
rect 4120 567208 67364 567236
rect 4120 567196 4126 567208
rect 67358 567196 67364 567208
rect 67416 567196 67422 567248
rect 1104 566800 68000 566896
rect 519948 566800 582820 566896
rect 1104 566256 68000 566352
rect 519948 566256 582820 566352
rect 1104 565712 68000 565808
rect 519948 565712 582820 565808
rect 1104 565168 68000 565264
rect 519948 565168 582820 565264
rect 1104 564624 68000 564720
rect 519948 564624 582820 564720
rect 520734 564340 520740 564392
rect 520792 564380 520798 564392
rect 580166 564380 580172 564392
rect 520792 564352 580172 564380
rect 520792 564340 520798 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 1104 564080 68000 564176
rect 519948 564080 582820 564176
rect 1104 563536 68000 563632
rect 519948 563536 582820 563632
rect 1104 562992 68000 563088
rect 519948 562992 582820 563088
rect 1104 562448 68000 562544
rect 519948 562448 582820 562544
rect 1104 561904 68000 562000
rect 519948 561904 582820 562000
rect 1104 561360 68000 561456
rect 519948 561360 582820 561456
rect 1104 560816 68000 560912
rect 519948 560816 582820 560912
rect 1104 560272 68000 560368
rect 519948 560272 582820 560368
rect 1104 559728 68000 559824
rect 519948 559728 582820 559824
rect 1104 559184 68000 559280
rect 519948 559184 582820 559280
rect 1104 558640 68000 558736
rect 519948 558640 582820 558736
rect 1104 558096 68000 558192
rect 519948 558096 582820 558192
rect 1104 557552 68000 557648
rect 519948 557552 582820 557648
rect 1104 557008 68000 557104
rect 519948 557008 582820 557104
rect 1104 556464 68000 556560
rect 519948 556464 582820 556560
rect 3418 556180 3424 556232
rect 3476 556220 3482 556232
rect 67358 556220 67364 556232
rect 3476 556192 67364 556220
rect 3476 556180 3482 556192
rect 67358 556180 67364 556192
rect 67416 556180 67422 556232
rect 1104 555920 68000 556016
rect 519948 555920 582820 556016
rect 1104 555376 68000 555472
rect 519948 555376 582820 555472
rect 1104 554832 68000 554928
rect 519948 554832 582820 554928
rect 1104 554288 68000 554384
rect 519948 554288 582820 554384
rect 1104 553744 68000 553840
rect 519948 553744 582820 553840
rect 1104 553200 68000 553296
rect 519948 553200 582820 553296
rect 1104 552656 68000 552752
rect 519948 552656 582820 552752
rect 1104 552112 68000 552208
rect 519948 552112 582820 552208
rect 521010 551964 521016 552016
rect 521068 552004 521074 552016
rect 579982 552004 579988 552016
rect 521068 551976 579988 552004
rect 521068 551964 521074 551976
rect 579982 551964 579988 551976
rect 580040 551964 580046 552016
rect 1104 551568 68000 551664
rect 519948 551568 582820 551664
rect 1104 551024 68000 551120
rect 519948 551024 582820 551120
rect 1104 550480 68000 550576
rect 519948 550480 582820 550576
rect 1104 549936 68000 550032
rect 519948 549936 582820 550032
rect 1104 549392 68000 549488
rect 519948 549392 582820 549488
rect 1104 548848 68000 548944
rect 519948 548848 582820 548944
rect 1104 548304 68000 548400
rect 519948 548304 582820 548400
rect 1104 547760 68000 547856
rect 519948 547760 582820 547856
rect 1104 547216 68000 547312
rect 519948 547216 582820 547312
rect 1104 546672 68000 546768
rect 519948 546672 582820 546768
rect 1104 546128 68000 546224
rect 519948 546128 582820 546224
rect 1104 545584 68000 545680
rect 519948 545584 582820 545680
rect 2958 545164 2964 545216
rect 3016 545204 3022 545216
rect 66622 545204 66628 545216
rect 3016 545176 66628 545204
rect 3016 545164 3022 545176
rect 66622 545164 66628 545176
rect 66680 545164 66686 545216
rect 1104 545040 68000 545136
rect 519948 545040 582820 545136
rect 1104 544496 68000 544592
rect 519948 544496 582820 544592
rect 1104 543952 68000 544048
rect 519948 543952 582820 544048
rect 1104 543408 68000 543504
rect 519948 543408 582820 543504
rect 1104 542864 68000 542960
rect 519948 542864 582820 542960
rect 1104 542320 68000 542416
rect 519948 542320 582820 542416
rect 1104 541776 68000 541872
rect 519948 541776 582820 541872
rect 1104 541232 68000 541328
rect 519948 541232 582820 541328
rect 1104 540688 68000 540784
rect 519948 540688 582820 540784
rect 1104 540144 68000 540240
rect 519948 540144 582820 540240
rect 1104 539600 68000 539696
rect 519948 539600 582820 539696
rect 1104 539056 68000 539152
rect 519948 539056 582820 539152
rect 1104 538512 68000 538608
rect 519948 538512 582820 538608
rect 520918 538160 520924 538212
rect 520976 538200 520982 538212
rect 580166 538200 580172 538212
rect 520976 538172 580172 538200
rect 520976 538160 520982 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 1104 537968 68000 538064
rect 519948 537968 582820 538064
rect 1104 537424 68000 537520
rect 519948 537424 582820 537520
rect 1104 536880 68000 536976
rect 519948 536880 582820 536976
rect 1104 536336 68000 536432
rect 519948 536336 582820 536432
rect 1104 535792 68000 535888
rect 519948 535792 582820 535888
rect 1104 535248 68000 535344
rect 519948 535248 582820 535344
rect 1104 534704 68000 534800
rect 519948 534704 582820 534800
rect 1104 534160 68000 534256
rect 519948 534160 582820 534256
rect 3418 534080 3424 534132
rect 3476 534120 3482 534132
rect 67358 534120 67364 534132
rect 3476 534092 67364 534120
rect 3476 534080 3482 534092
rect 67358 534080 67364 534092
rect 67416 534080 67422 534132
rect 1104 533616 68000 533712
rect 519948 533616 582820 533712
rect 1104 533072 68000 533168
rect 519948 533072 582820 533168
rect 1104 532528 68000 532624
rect 519948 532528 582820 532624
rect 1104 531984 68000 532080
rect 519948 531984 582820 532080
rect 1104 531440 68000 531536
rect 519948 531440 582820 531536
rect 1104 530896 68000 530992
rect 519948 530896 582820 530992
rect 1104 530352 68000 530448
rect 519948 530352 582820 530448
rect 1104 529808 68000 529904
rect 519948 529808 582820 529904
rect 1104 529264 68000 529360
rect 519948 529264 582820 529360
rect 1104 528720 68000 528816
rect 519948 528720 582820 528816
rect 1104 528176 68000 528272
rect 519948 528176 582820 528272
rect 1104 527632 68000 527728
rect 519948 527632 582820 527728
rect 1104 527088 68000 527184
rect 519948 527088 582820 527184
rect 1104 526544 68000 526640
rect 519948 526544 582820 526640
rect 1104 526000 68000 526096
rect 519948 526000 582820 526096
rect 520918 525716 520924 525768
rect 520976 525756 520982 525768
rect 579798 525756 579804 525768
rect 520976 525728 579804 525756
rect 520976 525716 520982 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 1104 525456 68000 525552
rect 519948 525456 582820 525552
rect 1104 524912 68000 525008
rect 519948 524912 582820 525008
rect 1104 524368 68000 524464
rect 519948 524368 582820 524464
rect 1104 523824 68000 523920
rect 519948 523824 582820 523920
rect 1104 523280 68000 523376
rect 519948 523280 582820 523376
rect 3418 522996 3424 523048
rect 3476 523036 3482 523048
rect 66438 523036 66444 523048
rect 3476 523008 66444 523036
rect 3476 522996 3482 523008
rect 66438 522996 66444 523008
rect 66496 522996 66502 523048
rect 1104 522736 68000 522832
rect 519948 522736 582820 522832
rect 1104 522192 68000 522288
rect 519948 522192 582820 522288
rect 1104 521648 68000 521744
rect 519948 521648 582820 521744
rect 1104 521104 68000 521200
rect 519948 521104 582820 521200
rect 1104 520560 68000 520656
rect 519948 520560 582820 520656
rect 1104 520016 68000 520112
rect 519948 520016 582820 520112
rect 1104 519472 68000 519568
rect 519948 519472 582820 519568
rect 1104 518928 68000 519024
rect 519948 518928 582820 519024
rect 1104 518384 68000 518480
rect 519948 518384 582820 518480
rect 1104 517840 68000 517936
rect 519948 517840 582820 517936
rect 1104 517296 68000 517392
rect 519948 517296 582820 517392
rect 1104 516752 68000 516848
rect 519948 516752 582820 516848
rect 1104 516208 68000 516304
rect 519948 516208 582820 516304
rect 1104 515664 68000 515760
rect 519948 515664 582820 515760
rect 1104 515120 68000 515216
rect 519948 515120 582820 515216
rect 1104 514576 68000 514672
rect 519948 514576 582820 514672
rect 1104 514032 68000 514128
rect 519948 514032 582820 514128
rect 1104 513488 68000 513584
rect 519948 513488 582820 513584
rect 1104 512944 68000 513040
rect 519948 512944 582820 513040
rect 1104 512400 68000 512496
rect 519948 512400 582820 512496
rect 3418 511980 3424 512032
rect 3476 512020 3482 512032
rect 67358 512020 67364 512032
rect 3476 511992 67364 512020
rect 3476 511980 3482 511992
rect 67358 511980 67364 511992
rect 67416 511980 67422 512032
rect 1104 511856 68000 511952
rect 519948 511856 582820 511952
rect 520918 511776 520924 511828
rect 520976 511816 520982 511828
rect 580166 511816 580172 511828
rect 520976 511788 580172 511816
rect 520976 511776 520982 511788
rect 580166 511776 580172 511788
rect 580224 511776 580230 511828
rect 1104 511312 68000 511408
rect 519948 511312 582820 511408
rect 1104 510768 68000 510864
rect 519948 510768 582820 510864
rect 1104 510224 68000 510320
rect 519948 510224 582820 510320
rect 1104 509680 68000 509776
rect 519948 509680 582820 509776
rect 1104 509136 68000 509232
rect 519948 509136 582820 509232
rect 1104 508592 68000 508688
rect 519948 508592 582820 508688
rect 1104 508048 68000 508144
rect 519948 508048 582820 508144
rect 1104 507504 68000 507600
rect 519948 507504 582820 507600
rect 1104 506960 68000 507056
rect 519948 506960 582820 507056
rect 1104 506416 68000 506512
rect 519948 506416 582820 506512
rect 1104 505872 68000 505968
rect 519948 505872 582820 505968
rect 1104 505328 68000 505424
rect 519948 505328 582820 505424
rect 1104 504784 68000 504880
rect 519948 504784 582820 504880
rect 1104 504240 68000 504336
rect 519948 504240 582820 504336
rect 1104 503696 68000 503792
rect 519948 503696 582820 503792
rect 1104 503152 68000 503248
rect 519948 503152 582820 503248
rect 1104 502608 68000 502704
rect 519948 502608 582820 502704
rect 1104 502064 68000 502160
rect 519948 502064 582820 502160
rect 1104 501520 68000 501616
rect 519948 501520 582820 501616
rect 3510 501100 3516 501152
rect 3568 501140 3574 501152
rect 67450 501140 67456 501152
rect 3568 501112 67456 501140
rect 3568 501100 3574 501112
rect 67450 501100 67456 501112
rect 67508 501100 67514 501152
rect 1104 500976 68000 501072
rect 519948 500976 582820 501072
rect 1104 500432 68000 500528
rect 519948 500432 582820 500528
rect 1104 499888 68000 499984
rect 519948 499888 582820 499984
rect 1104 499344 68000 499440
rect 519948 499344 582820 499440
rect 1104 498800 68000 498896
rect 519948 498800 582820 498896
rect 1104 498256 68000 498352
rect 519948 498256 582820 498352
rect 521010 498108 521016 498160
rect 521068 498148 521074 498160
rect 580166 498148 580172 498160
rect 521068 498120 580172 498148
rect 521068 498108 521074 498120
rect 580166 498108 580172 498120
rect 580224 498108 580230 498160
rect 1104 497712 68000 497808
rect 519948 497712 582820 497808
rect 1104 497168 68000 497264
rect 519948 497168 582820 497264
rect 1104 496624 68000 496720
rect 519948 496624 582820 496720
rect 1104 496080 68000 496176
rect 519948 496080 582820 496176
rect 1104 495536 68000 495632
rect 519948 495536 582820 495632
rect 1104 494992 68000 495088
rect 519948 494992 582820 495088
rect 1104 494448 68000 494544
rect 519948 494448 582820 494544
rect 1104 493904 68000 494000
rect 519948 493904 582820 494000
rect 1104 493360 68000 493456
rect 519948 493360 582820 493456
rect 1104 492816 68000 492912
rect 519948 492816 582820 492912
rect 1104 492272 68000 492368
rect 519948 492272 582820 492368
rect 1104 491728 68000 491824
rect 519948 491728 582820 491824
rect 1104 491184 68000 491280
rect 519948 491184 582820 491280
rect 1104 490640 68000 490736
rect 519948 490640 582820 490736
rect 1104 490096 68000 490192
rect 519948 490096 582820 490192
rect 3418 489880 3424 489932
rect 3476 489920 3482 489932
rect 67450 489920 67456 489932
rect 3476 489892 67456 489920
rect 3476 489880 3482 489892
rect 67450 489880 67456 489892
rect 67508 489880 67514 489932
rect 1104 489552 68000 489648
rect 519948 489552 582820 489648
rect 1104 489008 68000 489104
rect 519948 489008 582820 489104
rect 1104 488464 68000 488560
rect 519948 488464 582820 488560
rect 1104 487920 68000 488016
rect 519948 487920 582820 488016
rect 1104 487376 68000 487472
rect 519948 487376 582820 487472
rect 1104 486832 68000 486928
rect 519948 486832 582820 486928
rect 1104 486288 68000 486384
rect 519948 486288 582820 486384
rect 1104 485744 68000 485840
rect 519948 485744 582820 485840
rect 520918 485664 520924 485716
rect 520976 485704 520982 485716
rect 580166 485704 580172 485716
rect 520976 485676 580172 485704
rect 520976 485664 520982 485676
rect 580166 485664 580172 485676
rect 580224 485664 580230 485716
rect 1104 485200 68000 485296
rect 519948 485200 582820 485296
rect 1104 484656 68000 484752
rect 519948 484656 582820 484752
rect 1104 484112 68000 484208
rect 519948 484112 582820 484208
rect 1104 483568 68000 483664
rect 519948 483568 582820 483664
rect 1104 483024 68000 483120
rect 519948 483024 582820 483120
rect 1104 482480 68000 482576
rect 519948 482480 582820 482576
rect 1104 481936 68000 482032
rect 519948 481936 582820 482032
rect 1104 481392 68000 481488
rect 519948 481392 582820 481488
rect 1104 480848 68000 480944
rect 519948 480848 582820 480944
rect 1104 480304 68000 480400
rect 519948 480304 582820 480400
rect 1104 479760 68000 479856
rect 519948 479760 582820 479856
rect 1104 479216 68000 479312
rect 519948 479216 582820 479312
rect 3510 478864 3516 478916
rect 3568 478904 3574 478916
rect 67358 478904 67364 478916
rect 3568 478876 67364 478904
rect 3568 478864 3574 478876
rect 67358 478864 67364 478876
rect 67416 478864 67422 478916
rect 1104 478672 68000 478768
rect 519948 478672 582820 478768
rect 1104 478128 68000 478224
rect 519948 478128 582820 478224
rect 1104 477584 68000 477680
rect 519948 477584 582820 477680
rect 1104 477040 68000 477136
rect 519948 477040 582820 477136
rect 1104 476496 68000 476592
rect 519948 476496 582820 476592
rect 1104 475952 68000 476048
rect 519948 475952 582820 476048
rect 1104 475408 68000 475504
rect 519948 475408 582820 475504
rect 1104 474864 68000 474960
rect 519948 474864 582820 474960
rect 1104 474320 68000 474416
rect 519948 474320 582820 474416
rect 1104 473776 68000 473872
rect 519948 473776 582820 473872
rect 1104 473232 68000 473328
rect 519948 473232 582820 473328
rect 1104 472688 68000 472784
rect 519948 472688 582820 472784
rect 1104 472144 68000 472240
rect 519948 472144 582820 472240
rect 521010 471928 521016 471980
rect 521068 471968 521074 471980
rect 580166 471968 580172 471980
rect 521068 471940 580172 471968
rect 521068 471928 521074 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 1104 471600 68000 471696
rect 519948 471600 582820 471696
rect 1104 471056 68000 471152
rect 519948 471056 582820 471152
rect 1104 470512 68000 470608
rect 519948 470512 582820 470608
rect 1104 469968 68000 470064
rect 519948 469968 582820 470064
rect 1104 469424 68000 469520
rect 519948 469424 582820 469520
rect 1104 468880 68000 468976
rect 519948 468880 582820 468976
rect 1104 468336 68000 468432
rect 519948 468336 582820 468432
rect 1104 467792 68000 467888
rect 519948 467792 582820 467888
rect 1104 467248 68000 467344
rect 519948 467248 582820 467344
rect 1104 466704 68000 466800
rect 519948 466704 582820 466800
rect 3418 466420 3424 466472
rect 3476 466460 3482 466472
rect 66990 466460 66996 466472
rect 3476 466432 66996 466460
rect 3476 466420 3482 466432
rect 66990 466420 66996 466432
rect 67048 466420 67054 466472
rect 1104 466160 68000 466256
rect 519948 466160 582820 466256
rect 1104 465616 68000 465712
rect 519948 465616 582820 465712
rect 1104 465072 68000 465168
rect 519948 465072 582820 465168
rect 1104 464528 68000 464624
rect 519948 464528 582820 464624
rect 1104 463984 68000 464080
rect 519948 463984 582820 464080
rect 1104 463440 68000 463536
rect 519948 463440 582820 463536
rect 1104 462896 68000 462992
rect 519948 462896 582820 462992
rect 1104 462352 68000 462448
rect 519948 462352 582820 462448
rect 1104 461808 68000 461904
rect 519948 461808 582820 461904
rect 1104 461264 68000 461360
rect 519948 461264 582820 461360
rect 1104 460720 68000 460816
rect 519948 460720 582820 460816
rect 1104 460176 68000 460272
rect 519948 460176 582820 460272
rect 1104 459632 68000 459728
rect 519948 459632 582820 459728
rect 1104 459088 68000 459184
rect 519948 459088 582820 459184
rect 1104 458544 68000 458640
rect 519948 458544 582820 458640
rect 520918 458124 520924 458176
rect 520976 458164 520982 458176
rect 580166 458164 580172 458176
rect 520976 458136 580172 458164
rect 520976 458124 520982 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 1104 458000 68000 458096
rect 519948 458000 582820 458096
rect 1104 457456 68000 457552
rect 519948 457456 582820 457552
rect 1104 456912 68000 457008
rect 519948 456912 582820 457008
rect 1104 456368 68000 456464
rect 519948 456368 582820 456464
rect 1104 455824 68000 455920
rect 519948 455824 582820 455920
rect 3510 455404 3516 455456
rect 3568 455444 3574 455456
rect 67358 455444 67364 455456
rect 3568 455416 67364 455444
rect 3568 455404 3574 455416
rect 67358 455404 67364 455416
rect 67416 455404 67422 455456
rect 1104 455280 68000 455376
rect 519948 455280 582820 455376
rect 1104 454736 68000 454832
rect 519948 454736 582820 454832
rect 1104 454192 68000 454288
rect 519948 454192 582820 454288
rect 1104 453648 68000 453744
rect 519948 453648 582820 453744
rect 1104 453104 68000 453200
rect 519948 453104 582820 453200
rect 1104 452560 68000 452656
rect 519948 452560 582820 452656
rect 1104 452016 68000 452112
rect 519948 452016 582820 452112
rect 1104 451472 68000 451568
rect 519948 451472 582820 451568
rect 1104 450928 68000 451024
rect 519948 450928 582820 451024
rect 1104 450384 68000 450480
rect 519948 450384 582820 450480
rect 1104 449840 68000 449936
rect 519948 449840 582820 449936
rect 1104 449296 68000 449392
rect 519948 449296 582820 449392
rect 1104 448752 68000 448848
rect 519948 448752 582820 448848
rect 1104 448208 68000 448304
rect 519948 448208 582820 448304
rect 1104 447664 68000 447760
rect 519948 447664 582820 447760
rect 1104 447120 68000 447216
rect 519948 447120 582820 447216
rect 1104 446576 68000 446672
rect 519948 446576 582820 446672
rect 1104 446032 68000 446128
rect 519948 446032 582820 446128
rect 521102 445680 521108 445732
rect 521160 445720 521166 445732
rect 580166 445720 580172 445732
rect 521160 445692 580172 445720
rect 521160 445680 521166 445692
rect 580166 445680 580172 445692
rect 580224 445680 580230 445732
rect 1104 445488 68000 445584
rect 519948 445488 582820 445584
rect 1104 444944 68000 445040
rect 519948 444944 582820 445040
rect 3418 444524 3424 444576
rect 3476 444564 3482 444576
rect 66714 444564 66720 444576
rect 3476 444536 66720 444564
rect 3476 444524 3482 444536
rect 66714 444524 66720 444536
rect 66772 444524 66778 444576
rect 1104 444400 68000 444496
rect 519948 444400 582820 444496
rect 1104 443856 68000 443952
rect 519948 443856 582820 443952
rect 1104 443312 68000 443408
rect 519948 443312 582820 443408
rect 1104 442768 68000 442864
rect 519948 442768 582820 442864
rect 1104 442224 68000 442320
rect 519948 442224 582820 442320
rect 1104 441680 68000 441776
rect 519948 441680 582820 441776
rect 1104 441136 68000 441232
rect 519948 441136 582820 441232
rect 1104 440592 68000 440688
rect 519948 440592 582820 440688
rect 1104 440048 68000 440144
rect 519948 440048 582820 440144
rect 1104 439504 68000 439600
rect 519948 439504 582820 439600
rect 1104 438960 68000 439056
rect 519948 438960 582820 439056
rect 1104 438416 68000 438512
rect 519948 438416 582820 438512
rect 1104 437872 68000 437968
rect 519948 437872 582820 437968
rect 1104 437328 68000 437424
rect 519948 437328 582820 437424
rect 1104 436784 68000 436880
rect 519948 436784 582820 436880
rect 1104 436240 68000 436336
rect 519948 436240 582820 436336
rect 1104 435696 68000 435792
rect 519948 435696 582820 435792
rect 1104 435152 68000 435248
rect 519948 435152 582820 435248
rect 1104 434608 68000 434704
rect 519948 434608 582820 434704
rect 1104 434064 68000 434160
rect 519948 434064 582820 434160
rect 1104 433520 68000 433616
rect 519948 433520 582820 433616
rect 3602 433304 3608 433356
rect 3660 433344 3666 433356
rect 67174 433344 67180 433356
rect 3660 433316 67180 433344
rect 3660 433304 3666 433316
rect 67174 433304 67180 433316
rect 67232 433304 67238 433356
rect 1104 432976 68000 433072
rect 519948 432976 582820 433072
rect 1104 432432 68000 432528
rect 519948 432432 582820 432528
rect 1104 431888 68000 431984
rect 519948 431888 582820 431984
rect 521010 431808 521016 431860
rect 521068 431848 521074 431860
rect 580166 431848 580172 431860
rect 521068 431820 580172 431848
rect 521068 431808 521074 431820
rect 580166 431808 580172 431820
rect 580224 431808 580230 431860
rect 1104 431344 68000 431440
rect 519948 431344 582820 431440
rect 1104 430800 68000 430896
rect 519948 430800 582820 430896
rect 1104 430256 68000 430352
rect 519948 430256 582820 430352
rect 1104 429712 68000 429808
rect 519948 429712 582820 429808
rect 1104 429168 68000 429264
rect 519948 429168 582820 429264
rect 1104 428624 68000 428720
rect 519948 428624 582820 428720
rect 1104 428080 68000 428176
rect 519948 428080 582820 428176
rect 1104 427536 68000 427632
rect 519948 427536 582820 427632
rect 1104 426992 68000 427088
rect 519948 426992 582820 427088
rect 1104 426448 68000 426544
rect 519948 426448 582820 426544
rect 1104 425904 68000 426000
rect 519948 425904 582820 426000
rect 1104 425360 68000 425456
rect 519948 425360 582820 425456
rect 1104 424816 68000 424912
rect 519948 424816 582820 424912
rect 1104 424272 68000 424368
rect 519948 424272 582820 424368
rect 1104 423728 68000 423824
rect 519948 423728 582820 423824
rect 1104 423184 68000 423280
rect 519948 423184 582820 423280
rect 1104 422640 68000 422736
rect 519948 422640 582820 422736
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 66806 422328 66812 422340
rect 3568 422300 66812 422328
rect 3568 422288 3574 422300
rect 66806 422288 66812 422300
rect 66864 422288 66870 422340
rect 1104 422096 68000 422192
rect 519948 422096 582820 422192
rect 1104 421552 68000 421648
rect 519948 421552 582820 421648
rect 1104 421008 68000 421104
rect 519948 421008 582820 421104
rect 1104 420464 68000 420560
rect 519948 420464 582820 420560
rect 1104 419920 68000 420016
rect 519948 419920 582820 420016
rect 1104 419376 68000 419472
rect 519948 419376 582820 419472
rect 520918 419296 520924 419348
rect 520976 419336 520982 419348
rect 580166 419336 580172 419348
rect 520976 419308 580172 419336
rect 520976 419296 520982 419308
rect 580166 419296 580172 419308
rect 580224 419296 580230 419348
rect 1104 418832 68000 418928
rect 519948 418832 582820 418928
rect 1104 418288 68000 418384
rect 519948 418288 582820 418384
rect 1104 417744 68000 417840
rect 519948 417744 582820 417840
rect 1104 417200 68000 417296
rect 519948 417200 582820 417296
rect 1104 416656 68000 416752
rect 519948 416656 582820 416752
rect 1104 416112 68000 416208
rect 519948 416112 582820 416208
rect 1104 415568 68000 415664
rect 519948 415568 582820 415664
rect 1104 415024 68000 415120
rect 519948 415024 582820 415120
rect 1104 414480 68000 414576
rect 519948 414480 582820 414576
rect 1104 413936 68000 414032
rect 519948 413936 582820 414032
rect 1104 413392 68000 413488
rect 519948 413392 582820 413488
rect 1104 412848 68000 412944
rect 519948 412848 582820 412944
rect 1104 412304 68000 412400
rect 519948 412304 582820 412400
rect 1104 411760 68000 411856
rect 519948 411760 582820 411856
rect 3418 411340 3424 411392
rect 3476 411380 3482 411392
rect 67266 411380 67272 411392
rect 3476 411352 67272 411380
rect 3476 411340 3482 411352
rect 67266 411340 67272 411352
rect 67324 411340 67330 411392
rect 1104 411216 68000 411312
rect 519948 411216 582820 411312
rect 1104 410672 68000 410768
rect 519948 410672 582820 410768
rect 1104 410128 68000 410224
rect 519948 410128 582820 410224
rect 1104 409584 68000 409680
rect 519948 409584 582820 409680
rect 1104 409040 68000 409136
rect 519948 409040 582820 409136
rect 1104 408496 68000 408592
rect 519948 408496 582820 408592
rect 1104 407952 68000 408048
rect 519948 407952 582820 408048
rect 1104 407408 68000 407504
rect 519948 407408 582820 407504
rect 1104 406864 68000 406960
rect 519948 406864 582820 406960
rect 1104 406320 68000 406416
rect 519948 406320 582820 406416
rect 1104 405776 68000 405872
rect 519948 405776 582820 405872
rect 521010 405628 521016 405680
rect 521068 405668 521074 405680
rect 580166 405668 580172 405680
rect 521068 405640 580172 405668
rect 521068 405628 521074 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 1104 405232 68000 405328
rect 519948 405232 582820 405328
rect 1104 404688 68000 404784
rect 519948 404688 582820 404784
rect 1104 404144 68000 404240
rect 519948 404144 582820 404240
rect 1104 403600 68000 403696
rect 519948 403600 582820 403696
rect 1104 403056 68000 403152
rect 519948 403056 582820 403152
rect 1104 402512 68000 402608
rect 519948 402512 582820 402608
rect 1104 401968 68000 402064
rect 519948 401968 582820 402064
rect 1104 401424 68000 401520
rect 519948 401424 582820 401520
rect 1104 400880 68000 400976
rect 519948 400880 582820 400976
rect 1104 400336 68000 400432
rect 519948 400336 582820 400432
rect 3602 400188 3608 400240
rect 3660 400228 3666 400240
rect 67450 400228 67456 400240
rect 3660 400200 67456 400228
rect 3660 400188 3666 400200
rect 67450 400188 67456 400200
rect 67508 400188 67514 400240
rect 1104 399792 68000 399888
rect 519948 399792 582820 399888
rect 1104 399248 68000 399344
rect 519948 399248 582820 399344
rect 1104 398704 68000 398800
rect 519948 398704 582820 398800
rect 1104 398160 68000 398256
rect 519948 398160 582820 398256
rect 1104 397616 68000 397712
rect 519948 397616 582820 397712
rect 1104 397072 68000 397168
rect 519948 397072 582820 397168
rect 1104 396528 68000 396624
rect 519948 396528 582820 396624
rect 1104 395984 68000 396080
rect 519948 395984 582820 396080
rect 1104 395440 68000 395536
rect 519948 395440 582820 395536
rect 1104 394896 68000 394992
rect 519948 394896 582820 394992
rect 1104 394352 68000 394448
rect 519948 394352 582820 394448
rect 1104 393808 68000 393904
rect 519948 393808 582820 393904
rect 1104 393264 68000 393360
rect 519948 393264 582820 393360
rect 1104 392720 68000 392816
rect 519948 392720 582820 392816
rect 1104 392176 68000 392272
rect 519948 392176 582820 392272
rect 520918 391892 520924 391944
rect 520976 391932 520982 391944
rect 580166 391932 580172 391944
rect 520976 391904 580172 391932
rect 520976 391892 520982 391904
rect 580166 391892 580172 391904
rect 580224 391892 580230 391944
rect 1104 391632 68000 391728
rect 519948 391632 582820 391728
rect 1104 391088 68000 391184
rect 519948 391088 582820 391184
rect 1104 390544 68000 390640
rect 519948 390544 582820 390640
rect 1104 390000 68000 390096
rect 519948 390000 582820 390096
rect 1104 389456 68000 389552
rect 519948 389456 582820 389552
rect 3510 389172 3516 389224
rect 3568 389212 3574 389224
rect 67358 389212 67364 389224
rect 3568 389184 67364 389212
rect 3568 389172 3574 389184
rect 67358 389172 67364 389184
rect 67416 389172 67422 389224
rect 1104 388912 68000 389008
rect 519948 388912 582820 389008
rect 1104 388368 68000 388464
rect 519948 388368 582820 388464
rect 1104 387824 68000 387920
rect 519948 387824 582820 387920
rect 1104 387280 68000 387376
rect 519948 387280 582820 387376
rect 1104 386736 68000 386832
rect 519948 386736 582820 386832
rect 1104 386192 68000 386288
rect 519948 386192 582820 386288
rect 1104 385648 68000 385744
rect 519948 385648 582820 385744
rect 1104 385104 68000 385200
rect 519948 385104 582820 385200
rect 1104 384560 68000 384656
rect 519948 384560 582820 384656
rect 1104 384016 68000 384112
rect 519948 384016 582820 384112
rect 1104 383472 68000 383568
rect 519948 383472 582820 383568
rect 1104 382928 68000 383024
rect 519948 382928 582820 383024
rect 1104 382384 68000 382480
rect 519948 382384 582820 382480
rect 1104 381840 68000 381936
rect 519948 381840 582820 381936
rect 1104 381296 68000 381392
rect 519948 381296 582820 381392
rect 1104 380752 68000 380848
rect 519948 380752 582820 380848
rect 1104 380208 68000 380304
rect 519948 380208 582820 380304
rect 1104 379664 68000 379760
rect 519948 379664 582820 379760
rect 521102 379448 521108 379500
rect 521160 379488 521166 379500
rect 580166 379488 580172 379500
rect 521160 379460 580172 379488
rect 521160 379448 521166 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 1104 379120 68000 379216
rect 519948 379120 582820 379216
rect 1104 378576 68000 378672
rect 519948 378576 582820 378672
rect 3418 378156 3424 378208
rect 3476 378196 3482 378208
rect 67358 378196 67364 378208
rect 3476 378168 67364 378196
rect 3476 378156 3482 378168
rect 67358 378156 67364 378168
rect 67416 378156 67422 378208
rect 1104 378032 68000 378128
rect 519948 378032 582820 378128
rect 1104 377488 68000 377584
rect 519948 377488 582820 377584
rect 1104 376944 68000 377040
rect 519948 376944 582820 377040
rect 1104 376400 68000 376496
rect 519948 376400 582820 376496
rect 1104 375856 68000 375952
rect 519948 375856 582820 375952
rect 1104 375312 68000 375408
rect 519948 375312 582820 375408
rect 1104 374768 68000 374864
rect 519948 374768 582820 374864
rect 1104 374224 68000 374320
rect 519948 374224 582820 374320
rect 1104 373680 68000 373776
rect 519948 373680 582820 373776
rect 1104 373136 68000 373232
rect 519948 373136 582820 373232
rect 1104 372592 68000 372688
rect 519948 372592 582820 372688
rect 1104 372048 68000 372144
rect 519948 372048 582820 372144
rect 1104 371504 68000 371600
rect 519948 371504 582820 371600
rect 1104 370960 68000 371056
rect 519948 370960 582820 371056
rect 1104 370416 68000 370512
rect 519948 370416 582820 370512
rect 1104 369872 68000 369968
rect 519948 369872 582820 369968
rect 1104 369328 68000 369424
rect 519948 369328 582820 369424
rect 1104 368784 68000 368880
rect 519948 368784 582820 368880
rect 1104 368240 68000 368336
rect 519948 368240 582820 368336
rect 1104 367696 68000 367792
rect 519948 367696 582820 367792
rect 1104 367152 68000 367248
rect 519948 367152 582820 367248
rect 3694 367072 3700 367124
rect 3752 367112 3758 367124
rect 67358 367112 67364 367124
rect 3752 367084 67364 367112
rect 3752 367072 3758 367084
rect 67358 367072 67364 367084
rect 67416 367072 67422 367124
rect 1104 366608 68000 366704
rect 519948 366608 582820 366704
rect 1104 366064 68000 366160
rect 519948 366064 582820 366160
rect 521010 365644 521016 365696
rect 521068 365684 521074 365696
rect 580166 365684 580172 365696
rect 521068 365656 580172 365684
rect 521068 365644 521074 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 1104 365520 68000 365616
rect 519948 365520 582820 365616
rect 1104 364976 68000 365072
rect 519948 364976 582820 365072
rect 1104 364432 68000 364528
rect 519948 364432 582820 364528
rect 1104 363888 68000 363984
rect 519948 363888 582820 363984
rect 1104 363344 68000 363440
rect 519948 363344 582820 363440
rect 1104 362800 68000 362896
rect 519948 362800 582820 362896
rect 1104 362256 68000 362352
rect 519948 362256 582820 362352
rect 1104 361712 68000 361808
rect 519948 361712 582820 361808
rect 1104 361168 68000 361264
rect 519948 361168 582820 361264
rect 1104 360624 68000 360720
rect 519948 360624 582820 360720
rect 1104 360080 68000 360176
rect 519948 360080 582820 360176
rect 1104 359536 68000 359632
rect 519948 359536 582820 359632
rect 1104 358992 68000 359088
rect 519948 358992 582820 359088
rect 1104 358448 68000 358544
rect 519948 358448 582820 358544
rect 1104 357904 68000 358000
rect 519948 357904 582820 358000
rect 1104 357360 68000 357456
rect 519948 357360 582820 357456
rect 1104 356816 68000 356912
rect 519948 356816 582820 356912
rect 1104 356272 68000 356368
rect 519948 356272 582820 356368
rect 3602 356056 3608 356108
rect 3660 356096 3666 356108
rect 67358 356096 67364 356108
rect 3660 356068 67364 356096
rect 3660 356056 3666 356068
rect 67358 356056 67364 356068
rect 67416 356056 67422 356108
rect 1104 355728 68000 355824
rect 519948 355728 582820 355824
rect 1104 355184 68000 355280
rect 519948 355184 582820 355280
rect 1104 354640 68000 354736
rect 519948 354640 582820 354736
rect 1104 354096 68000 354192
rect 519948 354096 582820 354192
rect 1104 353552 68000 353648
rect 519948 353552 582820 353648
rect 520918 353200 520924 353252
rect 520976 353240 520982 353252
rect 580166 353240 580172 353252
rect 520976 353212 580172 353240
rect 520976 353200 520982 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 1104 353008 68000 353104
rect 519948 353008 582820 353104
rect 1104 352464 68000 352560
rect 519948 352464 582820 352560
rect 1104 351920 68000 352016
rect 519948 351920 582820 352016
rect 1104 351376 68000 351472
rect 519948 351376 582820 351472
rect 1104 350832 68000 350928
rect 519948 350832 582820 350928
rect 1104 350288 68000 350384
rect 519948 350288 582820 350384
rect 1104 349744 68000 349840
rect 519948 349744 582820 349840
rect 1104 349200 68000 349296
rect 519948 349200 582820 349296
rect 1104 348656 68000 348752
rect 519948 348656 582820 348752
rect 1104 348112 68000 348208
rect 519948 348112 582820 348208
rect 1104 347568 68000 347664
rect 519948 347568 582820 347664
rect 1104 347024 68000 347120
rect 519948 347024 582820 347120
rect 1104 346480 68000 346576
rect 519948 346480 582820 346576
rect 1104 345936 68000 346032
rect 519948 345936 582820 346032
rect 1104 345392 68000 345488
rect 519948 345392 582820 345488
rect 1104 344848 68000 344944
rect 519948 344848 582820 344944
rect 1104 344304 68000 344400
rect 519948 344304 582820 344400
rect 1104 343760 68000 343856
rect 519948 343760 582820 343856
rect 3510 343612 3516 343664
rect 3568 343652 3574 343664
rect 67358 343652 67364 343664
rect 3568 343624 67364 343652
rect 3568 343612 3574 343624
rect 67358 343612 67364 343624
rect 67416 343612 67422 343664
rect 1104 343216 68000 343312
rect 519948 343216 582820 343312
rect 1104 342672 68000 342768
rect 519948 342672 582820 342768
rect 1104 342128 68000 342224
rect 519948 342128 582820 342224
rect 1104 341584 68000 341680
rect 519948 341584 582820 341680
rect 1104 341040 68000 341136
rect 519948 341040 582820 341136
rect 1104 340496 68000 340592
rect 519948 340496 582820 340592
rect 1104 339952 68000 340048
rect 519948 339952 582820 340048
rect 1104 339408 68000 339504
rect 519948 339408 582820 339504
rect 521194 339328 521200 339380
rect 521252 339368 521258 339380
rect 580166 339368 580172 339380
rect 521252 339340 580172 339368
rect 521252 339328 521258 339340
rect 580166 339328 580172 339340
rect 580224 339328 580230 339380
rect 1104 338864 68000 338960
rect 519948 338864 582820 338960
rect 1104 338320 68000 338416
rect 519948 338320 582820 338416
rect 1104 337776 68000 337872
rect 519948 337776 582820 337872
rect 1104 337232 68000 337328
rect 519948 337232 582820 337328
rect 1104 336688 68000 336784
rect 519948 336688 582820 336784
rect 1104 336144 68000 336240
rect 519948 336144 582820 336240
rect 1104 335600 68000 335696
rect 519948 335600 582820 335696
rect 1104 335056 68000 335152
rect 519948 335056 582820 335152
rect 1104 334512 68000 334608
rect 519948 334512 582820 334608
rect 1104 333968 68000 334064
rect 519948 333968 582820 334064
rect 1104 333424 68000 333520
rect 519948 333424 582820 333520
rect 1104 332880 68000 332976
rect 519948 332880 582820 332976
rect 3418 332596 3424 332648
rect 3476 332636 3482 332648
rect 67174 332636 67180 332648
rect 3476 332608 67180 332636
rect 3476 332596 3482 332608
rect 67174 332596 67180 332608
rect 67232 332596 67238 332648
rect 1104 332336 68000 332432
rect 519948 332336 582820 332432
rect 1104 331792 68000 331888
rect 519948 331792 582820 331888
rect 1104 331248 68000 331344
rect 519948 331248 582820 331344
rect 1104 330704 68000 330800
rect 519948 330704 582820 330800
rect 1104 330160 68000 330256
rect 519948 330160 582820 330256
rect 1104 329616 68000 329712
rect 519948 329616 582820 329712
rect 1104 329072 68000 329168
rect 519948 329072 582820 329168
rect 1104 328528 68000 328624
rect 519948 328528 582820 328624
rect 1104 327984 68000 328080
rect 519948 327984 582820 328080
rect 1104 327440 68000 327536
rect 519948 327440 582820 327536
rect 1104 326896 68000 326992
rect 519948 326896 582820 326992
rect 1104 326352 68000 326448
rect 519948 326352 582820 326448
rect 1104 325808 68000 325904
rect 519948 325808 582820 325904
rect 521102 325592 521108 325644
rect 521160 325632 521166 325644
rect 580166 325632 580172 325644
rect 521160 325604 580172 325632
rect 521160 325592 521166 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 1104 325264 68000 325360
rect 519948 325264 582820 325360
rect 1104 324720 68000 324816
rect 519948 324720 582820 324816
rect 1104 324176 68000 324272
rect 519948 324176 582820 324272
rect 1104 323632 68000 323728
rect 519948 323632 582820 323728
rect 1104 323088 68000 323184
rect 519948 323088 582820 323184
rect 1104 322544 68000 322640
rect 519948 322544 582820 322640
rect 1104 322000 68000 322096
rect 519948 322000 582820 322096
rect 3694 321580 3700 321632
rect 3752 321620 3758 321632
rect 67358 321620 67364 321632
rect 3752 321592 67364 321620
rect 3752 321580 3758 321592
rect 67358 321580 67364 321592
rect 67416 321580 67422 321632
rect 1104 321456 68000 321552
rect 519948 321456 582820 321552
rect 1104 320912 68000 321008
rect 519948 320912 582820 321008
rect 1104 320368 68000 320464
rect 519948 320368 582820 320464
rect 1104 319824 68000 319920
rect 519948 319824 582820 319920
rect 1104 319280 68000 319376
rect 519948 319280 582820 319376
rect 1104 318736 68000 318832
rect 519948 318736 582820 318832
rect 1104 318192 68000 318288
rect 519948 318192 582820 318288
rect 1104 317648 68000 317744
rect 519948 317648 582820 317744
rect 1104 317104 68000 317200
rect 519948 317104 582820 317200
rect 1104 316560 68000 316656
rect 519948 316560 582820 316656
rect 1104 316016 68000 316112
rect 519948 316016 582820 316112
rect 1104 315472 68000 315568
rect 519948 315472 582820 315568
rect 1104 314928 68000 315024
rect 519948 314928 582820 315024
rect 1104 314384 68000 314480
rect 519948 314384 582820 314480
rect 1104 313840 68000 313936
rect 519948 313840 582820 313936
rect 1104 313296 68000 313392
rect 519948 313296 582820 313392
rect 521010 313216 521016 313268
rect 521068 313256 521074 313268
rect 580166 313256 580172 313268
rect 521068 313228 580172 313256
rect 521068 313216 521074 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 1104 312752 68000 312848
rect 519948 312752 582820 312848
rect 1104 312208 68000 312304
rect 519948 312208 582820 312304
rect 1104 311664 68000 311760
rect 519948 311664 582820 311760
rect 1104 311120 68000 311216
rect 519948 311120 582820 311216
rect 1104 310576 68000 310672
rect 519948 310576 582820 310672
rect 3602 310496 3608 310548
rect 3660 310536 3666 310548
rect 66714 310536 66720 310548
rect 3660 310508 66720 310536
rect 3660 310496 3666 310508
rect 66714 310496 66720 310508
rect 66772 310496 66778 310548
rect 1104 310032 68000 310128
rect 519948 310032 582820 310128
rect 1104 309488 68000 309584
rect 519948 309488 582820 309584
rect 1104 308944 68000 309040
rect 519948 308944 582820 309040
rect 1104 308400 68000 308496
rect 519948 308400 582820 308496
rect 1104 307856 68000 307952
rect 519948 307856 582820 307952
rect 1104 307312 68000 307408
rect 519948 307312 582820 307408
rect 1104 306768 68000 306864
rect 519948 306768 582820 306864
rect 1104 306224 68000 306320
rect 519948 306224 582820 306320
rect 1104 305680 68000 305776
rect 519948 305680 582820 305776
rect 1104 305136 68000 305232
rect 519948 305136 582820 305232
rect 1104 304592 68000 304688
rect 519948 304592 582820 304688
rect 1104 304048 68000 304144
rect 519948 304048 582820 304144
rect 1104 303504 68000 303600
rect 519948 303504 582820 303600
rect 1104 302960 68000 303056
rect 519948 302960 582820 303056
rect 1104 302416 68000 302512
rect 519948 302416 582820 302512
rect 1104 301872 68000 301968
rect 519948 301872 582820 301968
rect 1104 301328 68000 301424
rect 519948 301328 582820 301424
rect 1104 300784 68000 300880
rect 519948 300784 582820 300880
rect 1104 300240 68000 300336
rect 519948 300240 582820 300336
rect 1104 299696 68000 299792
rect 519948 299696 582820 299792
rect 3510 299480 3516 299532
rect 3568 299520 3574 299532
rect 67358 299520 67364 299532
rect 3568 299492 67364 299520
rect 3568 299480 3574 299492
rect 67358 299480 67364 299492
rect 67416 299480 67422 299532
rect 520918 299412 520924 299464
rect 520976 299452 520982 299464
rect 580166 299452 580172 299464
rect 520976 299424 580172 299452
rect 520976 299412 520982 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 1104 299152 68000 299248
rect 519948 299152 582820 299248
rect 1104 298608 68000 298704
rect 519948 298608 582820 298704
rect 1104 298064 68000 298160
rect 519948 298064 582820 298160
rect 1104 297520 68000 297616
rect 519948 297520 582820 297616
rect 1104 296976 68000 297072
rect 519948 296976 582820 297072
rect 1104 296432 68000 296528
rect 519948 296432 582820 296528
rect 1104 295888 68000 295984
rect 519948 295888 582820 295984
rect 1104 295344 68000 295440
rect 519948 295344 582820 295440
rect 1104 294800 68000 294896
rect 519948 294800 582820 294896
rect 1104 294256 68000 294352
rect 519948 294256 582820 294352
rect 1104 293712 68000 293808
rect 519948 293712 582820 293808
rect 1104 293168 68000 293264
rect 519948 293168 582820 293264
rect 1104 292624 68000 292720
rect 519948 292624 582820 292720
rect 1104 292080 68000 292176
rect 519948 292080 582820 292176
rect 1104 291536 68000 291632
rect 519948 291536 582820 291632
rect 1104 290992 68000 291088
rect 519948 290992 582820 291088
rect 1104 290448 68000 290544
rect 519948 290448 582820 290544
rect 1104 289904 68000 290000
rect 519948 289904 582820 290000
rect 1104 289360 68000 289456
rect 519948 289360 582820 289456
rect 1104 288816 68000 288912
rect 519948 288816 582820 288912
rect 3418 288396 3424 288448
rect 3476 288436 3482 288448
rect 66438 288436 66444 288448
rect 3476 288408 66444 288436
rect 3476 288396 3482 288408
rect 66438 288396 66444 288408
rect 66496 288396 66502 288448
rect 1104 288272 68000 288368
rect 519948 288272 582820 288368
rect 1104 287728 68000 287824
rect 519948 287728 582820 287824
rect 1104 287184 68000 287280
rect 519948 287184 582820 287280
rect 1104 286640 68000 286736
rect 519948 286640 582820 286736
rect 1104 286096 68000 286192
rect 519948 286096 582820 286192
rect 1104 285552 68000 285648
rect 519948 285552 582820 285648
rect 521194 285472 521200 285524
rect 521252 285512 521258 285524
rect 580166 285512 580172 285524
rect 521252 285484 580172 285512
rect 521252 285472 521258 285484
rect 580166 285472 580172 285484
rect 580224 285472 580230 285524
rect 1104 285008 68000 285104
rect 519948 285008 582820 285104
rect 1104 284464 68000 284560
rect 519948 284464 582820 284560
rect 1104 283920 68000 284016
rect 519948 283920 582820 284016
rect 1104 283376 68000 283472
rect 519948 283376 582820 283472
rect 1104 282832 68000 282928
rect 519948 282832 582820 282928
rect 1104 282288 68000 282384
rect 519948 282288 582820 282384
rect 1104 281744 68000 281840
rect 519948 281744 582820 281840
rect 1104 281200 68000 281296
rect 519948 281200 582820 281296
rect 1104 280656 68000 280752
rect 519948 280656 582820 280752
rect 1104 280112 68000 280208
rect 519948 280112 582820 280208
rect 1104 279568 68000 279664
rect 519948 279568 582820 279664
rect 1104 279024 68000 279120
rect 519948 279024 582820 279120
rect 1104 278480 68000 278576
rect 519948 278480 582820 278576
rect 1104 277936 68000 278032
rect 519948 277936 582820 278032
rect 3786 277516 3792 277568
rect 3844 277556 3850 277568
rect 67358 277556 67364 277568
rect 3844 277528 67364 277556
rect 3844 277516 3850 277528
rect 67358 277516 67364 277528
rect 67416 277516 67422 277568
rect 1104 277392 68000 277488
rect 519948 277392 582820 277488
rect 1104 276848 68000 276944
rect 519948 276848 582820 276944
rect 1104 276304 68000 276400
rect 519948 276304 582820 276400
rect 1104 275760 68000 275856
rect 519948 275760 582820 275856
rect 1104 275216 68000 275312
rect 519948 275216 582820 275312
rect 1104 274672 68000 274768
rect 519948 274672 582820 274768
rect 1104 274128 68000 274224
rect 519948 274128 582820 274224
rect 1104 273584 68000 273680
rect 519948 273584 582820 273680
rect 521102 273164 521108 273216
rect 521160 273204 521166 273216
rect 580166 273204 580172 273216
rect 521160 273176 580172 273204
rect 521160 273164 521166 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 1104 273040 68000 273136
rect 519948 273040 582820 273136
rect 1104 272496 68000 272592
rect 519948 272496 582820 272592
rect 1104 271952 68000 272048
rect 519948 271952 582820 272048
rect 1104 271408 68000 271504
rect 519948 271408 582820 271504
rect 1104 270864 68000 270960
rect 519948 270864 582820 270960
rect 1104 270320 68000 270416
rect 519948 270320 582820 270416
rect 1104 269776 68000 269872
rect 519948 269776 582820 269872
rect 1104 269232 68000 269328
rect 519948 269232 582820 269328
rect 1104 268688 68000 268784
rect 519948 268688 582820 268784
rect 1104 268144 68000 268240
rect 519948 268144 582820 268240
rect 1104 267600 68000 267696
rect 519948 267600 582820 267696
rect 1104 267056 68000 267152
rect 519948 267056 582820 267152
rect 1104 266512 68000 266608
rect 519948 266512 582820 266608
rect 3694 266364 3700 266416
rect 3752 266404 3758 266416
rect 67358 266404 67364 266416
rect 3752 266376 67364 266404
rect 3752 266364 3758 266376
rect 67358 266364 67364 266376
rect 67416 266364 67422 266416
rect 1104 265968 68000 266064
rect 519948 265968 582820 266064
rect 1104 265424 68000 265520
rect 519948 265424 582820 265520
rect 1104 264880 68000 264976
rect 519948 264880 582820 264976
rect 1104 264336 68000 264432
rect 519948 264336 582820 264432
rect 1104 263792 68000 263888
rect 519948 263792 582820 263888
rect 1104 263248 68000 263344
rect 519948 263248 582820 263344
rect 1104 262704 68000 262800
rect 519948 262704 582820 262800
rect 1104 262160 68000 262256
rect 519948 262160 582820 262256
rect 1104 261616 68000 261712
rect 519948 261616 582820 261712
rect 1104 261072 68000 261168
rect 519948 261072 582820 261168
rect 1104 260528 68000 260624
rect 519948 260528 582820 260624
rect 1104 259984 68000 260080
rect 519948 259984 582820 260080
rect 1104 259440 68000 259536
rect 519948 259440 582820 259536
rect 521010 259360 521016 259412
rect 521068 259400 521074 259412
rect 580166 259400 580172 259412
rect 521068 259372 580172 259400
rect 521068 259360 521074 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 1104 258896 68000 258992
rect 519948 258896 582820 258992
rect 1104 258352 68000 258448
rect 519948 258352 582820 258448
rect 1104 257808 68000 257904
rect 519948 257808 582820 257904
rect 1104 257264 68000 257360
rect 519948 257264 582820 257360
rect 1104 256720 68000 256816
rect 519948 256720 582820 256816
rect 1104 256176 68000 256272
rect 519948 256176 582820 256272
rect 1104 255632 68000 255728
rect 519948 255632 582820 255728
rect 3602 255280 3608 255332
rect 3660 255320 3666 255332
rect 67358 255320 67364 255332
rect 3660 255292 67364 255320
rect 3660 255280 3666 255292
rect 67358 255280 67364 255292
rect 67416 255280 67422 255332
rect 1104 255088 68000 255184
rect 519948 255088 582820 255184
rect 1104 254544 68000 254640
rect 519948 254544 582820 254640
rect 1104 254000 68000 254096
rect 519948 254000 582820 254096
rect 1104 253456 68000 253552
rect 519948 253456 582820 253552
rect 1104 252912 68000 253008
rect 519948 252912 582820 253008
rect 1104 252368 68000 252464
rect 519948 252368 582820 252464
rect 1104 251824 68000 251920
rect 519948 251824 582820 251920
rect 1104 251280 68000 251376
rect 519948 251280 582820 251376
rect 1104 250736 68000 250832
rect 519948 250736 582820 250832
rect 1104 250192 68000 250288
rect 519948 250192 582820 250288
rect 1104 249648 68000 249744
rect 519948 249648 582820 249744
rect 1104 249104 68000 249200
rect 519948 249104 582820 249200
rect 1104 248560 68000 248656
rect 519948 248560 582820 248656
rect 1104 248016 68000 248112
rect 519948 248016 582820 248112
rect 1104 247472 68000 247568
rect 519948 247472 582820 247568
rect 1104 246928 68000 247024
rect 519948 246928 582820 247024
rect 1104 246384 68000 246480
rect 519948 246384 582820 246480
rect 1104 245840 68000 245936
rect 519948 245840 582820 245936
rect 520918 245556 520924 245608
rect 520976 245596 520982 245608
rect 580166 245596 580172 245608
rect 520976 245568 580172 245596
rect 520976 245556 520982 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 1104 245296 68000 245392
rect 519948 245296 582820 245392
rect 1104 244752 68000 244848
rect 519948 244752 582820 244848
rect 3510 244332 3516 244384
rect 3568 244372 3574 244384
rect 67358 244372 67364 244384
rect 3568 244344 67364 244372
rect 3568 244332 3574 244344
rect 67358 244332 67364 244344
rect 67416 244332 67422 244384
rect 1104 244208 68000 244304
rect 519948 244208 582820 244304
rect 1104 243664 68000 243760
rect 519948 243664 582820 243760
rect 1104 243120 68000 243216
rect 519948 243120 582820 243216
rect 1104 242576 68000 242672
rect 519948 242576 582820 242672
rect 1104 242032 68000 242128
rect 519948 242032 582820 242128
rect 1104 241488 68000 241584
rect 519948 241488 582820 241584
rect 1104 240944 68000 241040
rect 519948 240944 582820 241040
rect 1104 240400 68000 240496
rect 519948 240400 582820 240496
rect 1104 239856 68000 239952
rect 519948 239856 582820 239952
rect 1104 239312 68000 239408
rect 519948 239312 582820 239408
rect 1104 238768 68000 238864
rect 519948 238768 582820 238864
rect 1104 238224 68000 238320
rect 519948 238224 582820 238320
rect 1104 237680 68000 237776
rect 519948 237680 582820 237776
rect 1104 237136 68000 237232
rect 519948 237136 582820 237232
rect 1104 236592 68000 236688
rect 519948 236592 582820 236688
rect 1104 236048 68000 236144
rect 519948 236048 582820 236144
rect 1104 235504 68000 235600
rect 519948 235504 582820 235600
rect 1104 234960 68000 235056
rect 519948 234960 582820 235056
rect 1104 234416 68000 234512
rect 519948 234416 582820 234512
rect 1104 233872 68000 233968
rect 519948 233872 582820 233968
rect 1104 233328 68000 233424
rect 519948 233328 582820 233424
rect 3418 233248 3424 233300
rect 3476 233288 3482 233300
rect 67174 233288 67180 233300
rect 3476 233260 67180 233288
rect 3476 233248 3482 233260
rect 67174 233248 67180 233260
rect 67232 233248 67238 233300
rect 521286 233180 521292 233232
rect 521344 233220 521350 233232
rect 579982 233220 579988 233232
rect 521344 233192 579988 233220
rect 521344 233180 521350 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 1104 232784 68000 232880
rect 519948 232784 582820 232880
rect 1104 232240 68000 232336
rect 519948 232240 582820 232336
rect 1104 231696 68000 231792
rect 519948 231696 582820 231792
rect 1104 231152 68000 231248
rect 519948 231152 582820 231248
rect 1104 230608 68000 230704
rect 519948 230608 582820 230704
rect 1104 230064 68000 230160
rect 519948 230064 582820 230160
rect 1104 229520 68000 229616
rect 519948 229520 582820 229616
rect 1104 228976 68000 229072
rect 519948 228976 582820 229072
rect 1104 228432 68000 228528
rect 519948 228432 582820 228528
rect 1104 227888 68000 227984
rect 519948 227888 582820 227984
rect 1104 227344 68000 227440
rect 519948 227344 582820 227440
rect 1104 226800 68000 226896
rect 519948 226800 582820 226896
rect 1104 226256 68000 226352
rect 519948 226256 582820 226352
rect 1104 225712 68000 225808
rect 519948 225712 582820 225808
rect 1104 225168 68000 225264
rect 519948 225168 582820 225264
rect 1104 224624 68000 224720
rect 519948 224624 582820 224720
rect 1104 224080 68000 224176
rect 519948 224080 582820 224176
rect 1104 223536 68000 223632
rect 519948 223536 582820 223632
rect 1104 222992 68000 223088
rect 519948 222992 582820 223088
rect 1104 222448 68000 222544
rect 519948 222448 582820 222544
rect 1104 221904 68000 222000
rect 519948 221904 582820 222000
rect 1104 221360 68000 221456
rect 519948 221360 582820 221456
rect 3878 220940 3884 220992
rect 3936 220980 3942 220992
rect 67358 220980 67364 220992
rect 3936 220952 67364 220980
rect 3936 220940 3942 220952
rect 67358 220940 67364 220952
rect 67416 220940 67422 220992
rect 1104 220816 68000 220912
rect 519948 220816 582820 220912
rect 1104 220272 68000 220368
rect 519948 220272 582820 220368
rect 1104 219728 68000 219824
rect 519948 219728 582820 219824
rect 521194 219376 521200 219428
rect 521252 219416 521258 219428
rect 580166 219416 580172 219428
rect 521252 219388 580172 219416
rect 521252 219376 521258 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 1104 219184 68000 219280
rect 519948 219184 582820 219280
rect 1104 218640 68000 218736
rect 519948 218640 582820 218736
rect 1104 218096 68000 218192
rect 519948 218096 582820 218192
rect 1104 217552 68000 217648
rect 519948 217552 582820 217648
rect 1104 217008 68000 217104
rect 519948 217008 582820 217104
rect 1104 216464 68000 216560
rect 519948 216464 582820 216560
rect 1104 215920 68000 216016
rect 519948 215920 582820 216016
rect 1104 215376 68000 215472
rect 519948 215376 582820 215472
rect 1104 214832 68000 214928
rect 519948 214832 582820 214928
rect 1104 214288 68000 214384
rect 519948 214288 582820 214384
rect 1104 213744 68000 213840
rect 519948 213744 582820 213840
rect 1104 213200 68000 213296
rect 519948 213200 582820 213296
rect 1104 212656 68000 212752
rect 519948 212656 582820 212752
rect 1104 212112 68000 212208
rect 519948 212112 582820 212208
rect 1104 211568 68000 211664
rect 519948 211568 582820 211664
rect 1104 211024 68000 211120
rect 519948 211024 582820 211120
rect 1104 210480 68000 210576
rect 519948 210480 582820 210576
rect 1104 209936 68000 210032
rect 519948 209936 582820 210032
rect 3786 209788 3792 209840
rect 3844 209828 3850 209840
rect 67358 209828 67364 209840
rect 3844 209800 67364 209828
rect 3844 209788 3850 209800
rect 67358 209788 67364 209800
rect 67416 209788 67422 209840
rect 1104 209392 68000 209488
rect 519948 209392 582820 209488
rect 1104 208848 68000 208944
rect 519948 208848 582820 208944
rect 1104 208304 68000 208400
rect 519948 208304 582820 208400
rect 1104 207760 68000 207856
rect 519948 207760 582820 207856
rect 1104 207216 68000 207312
rect 519948 207216 582820 207312
rect 521102 206932 521108 206984
rect 521160 206972 521166 206984
rect 579798 206972 579804 206984
rect 521160 206944 579804 206972
rect 521160 206932 521166 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 1104 206672 68000 206768
rect 519948 206672 582820 206768
rect 1104 206128 68000 206224
rect 519948 206128 582820 206224
rect 1104 205584 68000 205680
rect 519948 205584 582820 205680
rect 1104 205040 68000 205136
rect 519948 205040 582820 205136
rect 1104 204496 68000 204592
rect 519948 204496 582820 204592
rect 1104 203952 68000 204048
rect 519948 203952 582820 204048
rect 1104 203408 68000 203504
rect 519948 203408 582820 203504
rect 1104 202864 68000 202960
rect 519948 202864 582820 202960
rect 1104 202320 68000 202416
rect 519948 202320 582820 202416
rect 1104 201776 68000 201872
rect 519948 201776 582820 201872
rect 1104 201232 68000 201328
rect 519948 201232 582820 201328
rect 1104 200688 68000 200784
rect 519948 200688 582820 200784
rect 1104 200144 68000 200240
rect 519948 200144 582820 200240
rect 1104 199600 68000 199696
rect 519948 199600 582820 199696
rect 1104 199056 68000 199152
rect 519948 199056 582820 199152
rect 3694 198704 3700 198756
rect 3752 198744 3758 198756
rect 67358 198744 67364 198756
rect 3752 198716 67364 198744
rect 3752 198704 3758 198716
rect 67358 198704 67364 198716
rect 67416 198704 67422 198756
rect 1104 198512 68000 198608
rect 519948 198512 582820 198608
rect 1104 197968 68000 198064
rect 519948 197968 582820 198064
rect 1104 197424 68000 197520
rect 519948 197424 582820 197520
rect 1104 196880 68000 196976
rect 519948 196880 582820 196976
rect 1104 196336 68000 196432
rect 519948 196336 582820 196432
rect 1104 195792 68000 195888
rect 519948 195792 582820 195888
rect 1104 195248 68000 195344
rect 519948 195248 582820 195344
rect 1104 194704 68000 194800
rect 519948 194704 582820 194800
rect 1104 194160 68000 194256
rect 519948 194160 582820 194256
rect 1104 193616 68000 193712
rect 519948 193616 582820 193712
rect 1104 193072 68000 193168
rect 519948 193072 582820 193168
rect 521010 192992 521016 193044
rect 521068 193032 521074 193044
rect 580166 193032 580172 193044
rect 521068 193004 580172 193032
rect 521068 192992 521074 193004
rect 580166 192992 580172 193004
rect 580224 192992 580230 193044
rect 1104 192528 68000 192624
rect 519948 192528 582820 192624
rect 1104 191984 68000 192080
rect 519948 191984 582820 192080
rect 1104 191440 68000 191536
rect 519948 191440 582820 191536
rect 1104 190896 68000 190992
rect 519948 190896 582820 190992
rect 1104 190352 68000 190448
rect 519948 190352 582820 190448
rect 1104 189808 68000 189904
rect 519948 189808 582820 189904
rect 1104 189264 68000 189360
rect 519948 189264 582820 189360
rect 1104 188720 68000 188816
rect 519948 188720 582820 188816
rect 1104 188176 68000 188272
rect 519948 188176 582820 188272
rect 3602 187756 3608 187808
rect 3660 187796 3666 187808
rect 67450 187796 67456 187808
rect 3660 187768 67456 187796
rect 3660 187756 3666 187768
rect 67450 187756 67456 187768
rect 67508 187756 67514 187808
rect 1104 187632 68000 187728
rect 519948 187632 582820 187728
rect 1104 187088 68000 187184
rect 519948 187088 582820 187184
rect 1104 186544 68000 186640
rect 519948 186544 582820 186640
rect 1104 186000 68000 186096
rect 519948 186000 582820 186096
rect 1104 185456 68000 185552
rect 519948 185456 582820 185552
rect 1104 184912 68000 185008
rect 519948 184912 582820 185008
rect 1104 184368 68000 184464
rect 519948 184368 582820 184464
rect 1104 183824 68000 183920
rect 519948 183824 582820 183920
rect 1104 183280 68000 183376
rect 519948 183280 582820 183376
rect 1104 182736 68000 182832
rect 519948 182736 582820 182832
rect 1104 182192 68000 182288
rect 519948 182192 582820 182288
rect 1104 181648 68000 181744
rect 519948 181648 582820 181744
rect 1104 181104 68000 181200
rect 519948 181104 582820 181200
rect 1104 180560 68000 180656
rect 519948 180560 582820 180656
rect 1104 180016 68000 180112
rect 519948 180016 582820 180112
rect 1104 179472 68000 179568
rect 519948 179472 582820 179568
rect 520918 179324 520924 179376
rect 520976 179364 520982 179376
rect 580166 179364 580172 179376
rect 520976 179336 580172 179364
rect 520976 179324 520982 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 1104 178928 68000 179024
rect 519948 178928 582820 179024
rect 1104 178384 68000 178480
rect 519948 178384 582820 178480
rect 1104 177840 68000 177936
rect 519948 177840 582820 177936
rect 1104 177296 68000 177392
rect 519948 177296 582820 177392
rect 1104 176752 68000 176848
rect 519948 176752 582820 176848
rect 3510 176672 3516 176724
rect 3568 176712 3574 176724
rect 67358 176712 67364 176724
rect 3568 176684 67364 176712
rect 3568 176672 3574 176684
rect 67358 176672 67364 176684
rect 67416 176672 67422 176724
rect 1104 176208 68000 176304
rect 519948 176208 582820 176304
rect 1104 175664 68000 175760
rect 519948 175664 582820 175760
rect 1104 175120 68000 175216
rect 519948 175120 582820 175216
rect 1104 174576 68000 174672
rect 519948 174576 582820 174672
rect 1104 174032 68000 174128
rect 519948 174032 582820 174128
rect 1104 173488 68000 173584
rect 519948 173488 582820 173584
rect 1104 172944 68000 173040
rect 519948 172944 582820 173040
rect 1104 172400 68000 172496
rect 519948 172400 582820 172496
rect 1104 171856 68000 171952
rect 519948 171856 582820 171952
rect 1104 171312 68000 171408
rect 519948 171312 582820 171408
rect 1104 170768 68000 170864
rect 519948 170768 582820 170864
rect 1104 170224 68000 170320
rect 519948 170224 582820 170320
rect 1104 169680 68000 169776
rect 519948 169680 582820 169776
rect 1104 169136 68000 169232
rect 519948 169136 582820 169232
rect 1104 168592 68000 168688
rect 519948 168592 582820 168688
rect 1104 168048 68000 168144
rect 519948 168048 582820 168144
rect 1104 167504 68000 167600
rect 519948 167504 582820 167600
rect 1104 166960 68000 167056
rect 519948 166960 582820 167056
rect 521378 166880 521384 166932
rect 521436 166920 521442 166932
rect 580166 166920 580172 166932
rect 521436 166892 580172 166920
rect 521436 166880 521442 166892
rect 580166 166880 580172 166892
rect 580224 166880 580230 166932
rect 1104 166416 68000 166512
rect 519948 166416 582820 166512
rect 1104 165872 68000 165968
rect 519948 165872 582820 165968
rect 3418 165588 3424 165640
rect 3476 165628 3482 165640
rect 67358 165628 67364 165640
rect 3476 165600 67364 165628
rect 3476 165588 3482 165600
rect 67358 165588 67364 165600
rect 67416 165588 67422 165640
rect 1104 165328 68000 165424
rect 519948 165328 582820 165424
rect 1104 164784 68000 164880
rect 519948 164784 582820 164880
rect 1104 164240 68000 164336
rect 519948 164240 582820 164336
rect 1104 163696 68000 163792
rect 519948 163696 582820 163792
rect 1104 163152 68000 163248
rect 519948 163152 582820 163248
rect 1104 162608 68000 162704
rect 519948 162608 582820 162704
rect 1104 162064 68000 162160
rect 519948 162064 582820 162160
rect 1104 161520 68000 161616
rect 519948 161520 582820 161616
rect 1104 160976 68000 161072
rect 519948 160976 582820 161072
rect 1104 160432 68000 160528
rect 519948 160432 582820 160528
rect 1104 159888 68000 159984
rect 519948 159888 582820 159984
rect 1104 159344 68000 159440
rect 519948 159344 582820 159440
rect 1104 158800 68000 158896
rect 519948 158800 582820 158896
rect 1104 158256 68000 158352
rect 519948 158256 582820 158352
rect 1104 157712 68000 157808
rect 519948 157712 582820 157808
rect 1104 157168 68000 157264
rect 519948 157168 582820 157264
rect 1104 156624 68000 156720
rect 519948 156624 582820 156720
rect 1104 156080 68000 156176
rect 519948 156080 582820 156176
rect 1104 155536 68000 155632
rect 519948 155536 582820 155632
rect 1104 154992 68000 155088
rect 519948 154992 582820 155088
rect 3970 154572 3976 154624
rect 4028 154612 4034 154624
rect 67266 154612 67272 154624
rect 4028 154584 67272 154612
rect 4028 154572 4034 154584
rect 67266 154572 67272 154584
rect 67324 154572 67330 154624
rect 1104 154448 68000 154544
rect 519948 154448 582820 154544
rect 1104 153904 68000 154000
rect 519948 153904 582820 154000
rect 1104 153360 68000 153456
rect 519948 153360 582820 153456
rect 521286 153144 521292 153196
rect 521344 153184 521350 153196
rect 580166 153184 580172 153196
rect 521344 153156 580172 153184
rect 521344 153144 521350 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 1104 152816 68000 152912
rect 519948 152816 582820 152912
rect 1104 152272 68000 152368
rect 519948 152272 582820 152368
rect 1104 151728 68000 151824
rect 519948 151728 582820 151824
rect 1104 151184 68000 151280
rect 519948 151184 582820 151280
rect 1104 150640 68000 150736
rect 519948 150640 582820 150736
rect 1104 150096 68000 150192
rect 519948 150096 582820 150192
rect 1104 149552 68000 149648
rect 519948 149552 582820 149648
rect 1104 149008 68000 149104
rect 519948 149008 582820 149104
rect 1104 148464 68000 148560
rect 519948 148464 582820 148560
rect 1104 147920 68000 148016
rect 519948 147920 582820 148016
rect 1104 147376 68000 147472
rect 519948 147376 582820 147472
rect 1104 146832 68000 146928
rect 519948 146832 582820 146928
rect 1104 146288 68000 146384
rect 519948 146288 582820 146384
rect 1104 145744 68000 145840
rect 519948 145744 582820 145840
rect 1104 145200 68000 145296
rect 519948 145200 582820 145296
rect 1104 144656 68000 144752
rect 519948 144656 582820 144752
rect 1104 144112 68000 144208
rect 519948 144112 582820 144208
rect 3878 143692 3884 143744
rect 3936 143732 3942 143744
rect 67358 143732 67364 143744
rect 3936 143704 67364 143732
rect 3936 143692 3942 143704
rect 67358 143692 67364 143704
rect 67416 143692 67422 143744
rect 1104 143568 68000 143664
rect 519948 143568 582820 143664
rect 1104 143024 68000 143120
rect 519948 143024 582820 143120
rect 1104 142480 68000 142576
rect 519948 142480 582820 142576
rect 1104 141936 68000 142032
rect 519948 141936 582820 142032
rect 1104 141392 68000 141488
rect 519948 141392 582820 141488
rect 1104 140848 68000 140944
rect 519948 140848 582820 140944
rect 1104 140304 68000 140400
rect 519948 140304 582820 140400
rect 1104 139760 68000 139856
rect 519948 139760 582820 139856
rect 521194 139340 521200 139392
rect 521252 139380 521258 139392
rect 580166 139380 580172 139392
rect 521252 139352 580172 139380
rect 521252 139340 521258 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 1104 139216 68000 139312
rect 519948 139216 582820 139312
rect 1104 138672 68000 138768
rect 519948 138672 582820 138768
rect 1104 138128 68000 138224
rect 519948 138128 582820 138224
rect 1104 137584 68000 137680
rect 519948 137584 582820 137680
rect 1104 137040 68000 137136
rect 519948 137040 582820 137136
rect 1104 136496 68000 136592
rect 519948 136496 582820 136592
rect 1104 135952 68000 136048
rect 519948 135952 582820 136048
rect 1104 135408 68000 135504
rect 519948 135408 582820 135504
rect 1104 134864 68000 134960
rect 519948 134864 582820 134960
rect 1104 134320 68000 134416
rect 519948 134320 582820 134416
rect 1104 133776 68000 133872
rect 519948 133776 582820 133872
rect 1104 133232 68000 133328
rect 519948 133232 582820 133328
rect 1104 132688 68000 132784
rect 519948 132688 582820 132784
rect 3786 132472 3792 132524
rect 3844 132512 3850 132524
rect 67174 132512 67180 132524
rect 3844 132484 67180 132512
rect 3844 132472 3850 132484
rect 67174 132472 67180 132484
rect 67232 132472 67238 132524
rect 1104 132144 68000 132240
rect 519948 132144 582820 132240
rect 1104 131600 68000 131696
rect 519948 131600 582820 131696
rect 1104 131056 68000 131152
rect 519948 131056 582820 131152
rect 1104 130512 68000 130608
rect 519948 130512 582820 130608
rect 1104 129968 68000 130064
rect 519948 129968 582820 130064
rect 1104 129424 68000 129520
rect 519948 129424 582820 129520
rect 1104 128880 68000 128976
rect 519948 128880 582820 128976
rect 1104 128336 68000 128432
rect 519948 128336 582820 128432
rect 1104 127792 68000 127888
rect 519948 127792 582820 127888
rect 1104 127248 68000 127344
rect 519948 127248 582820 127344
rect 521102 126896 521108 126948
rect 521160 126936 521166 126948
rect 580166 126936 580172 126948
rect 521160 126908 580172 126936
rect 521160 126896 521166 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 1104 126704 68000 126800
rect 519948 126704 582820 126800
rect 1104 126160 68000 126256
rect 519948 126160 582820 126256
rect 1104 125616 68000 125712
rect 519948 125616 582820 125712
rect 1104 125072 68000 125168
rect 519948 125072 582820 125168
rect 1104 124528 68000 124624
rect 519948 124528 582820 124624
rect 1104 123984 68000 124080
rect 519948 123984 582820 124080
rect 1104 123440 68000 123536
rect 519948 123440 582820 123536
rect 1104 122896 68000 122992
rect 519948 122896 582820 122992
rect 1104 122352 68000 122448
rect 519948 122352 582820 122448
rect 1104 121808 68000 121904
rect 519948 121808 582820 121904
rect 3694 121456 3700 121508
rect 3752 121496 3758 121508
rect 67358 121496 67364 121508
rect 3752 121468 67364 121496
rect 3752 121456 3758 121468
rect 67358 121456 67364 121468
rect 67416 121456 67422 121508
rect 1104 121264 68000 121360
rect 519948 121264 582820 121360
rect 1104 120720 68000 120816
rect 519948 120720 582820 120816
rect 1104 120176 68000 120272
rect 519948 120176 582820 120272
rect 1104 119632 68000 119728
rect 519948 119632 582820 119728
rect 1104 119088 68000 119184
rect 519948 119088 582820 119184
rect 1104 118544 68000 118640
rect 519948 118544 582820 118640
rect 1104 118000 68000 118096
rect 519948 118000 582820 118096
rect 1104 117456 68000 117552
rect 519948 117456 582820 117552
rect 1104 116912 68000 117008
rect 519948 116912 582820 117008
rect 1104 116368 68000 116464
rect 519948 116368 582820 116464
rect 1104 115824 68000 115920
rect 519948 115824 582820 115920
rect 1104 115280 68000 115376
rect 519948 115280 582820 115376
rect 1104 114736 68000 114832
rect 519948 114736 582820 114832
rect 1104 114192 68000 114288
rect 519948 114192 582820 114288
rect 1104 113648 68000 113744
rect 519948 113648 582820 113744
rect 1104 113104 68000 113200
rect 519948 113104 582820 113200
rect 521010 113024 521016 113076
rect 521068 113064 521074 113076
rect 580166 113064 580172 113076
rect 521068 113036 580172 113064
rect 521068 113024 521074 113036
rect 580166 113024 580172 113036
rect 580224 113024 580230 113076
rect 1104 112560 68000 112656
rect 519948 112560 582820 112656
rect 1104 112016 68000 112112
rect 519948 112016 582820 112112
rect 1104 111472 68000 111568
rect 519948 111472 582820 111568
rect 1104 110928 68000 111024
rect 519948 110928 582820 111024
rect 1104 110384 68000 110480
rect 519948 110384 582820 110480
rect 1104 109840 68000 109936
rect 519948 109840 582820 109936
rect 1104 109296 68000 109392
rect 519948 109296 582820 109392
rect 3602 109012 3608 109064
rect 3660 109052 3666 109064
rect 67358 109052 67364 109064
rect 3660 109024 67364 109052
rect 3660 109012 3666 109024
rect 67358 109012 67364 109024
rect 67416 109012 67422 109064
rect 1104 108752 68000 108848
rect 519948 108752 582820 108848
rect 1104 108208 68000 108304
rect 519948 108208 582820 108304
rect 1104 107664 68000 107760
rect 519948 107664 582820 107760
rect 1104 107120 68000 107216
rect 519948 107120 582820 107216
rect 1104 106576 68000 106672
rect 519948 106576 582820 106672
rect 1104 106032 68000 106128
rect 519948 106032 582820 106128
rect 1104 105488 68000 105584
rect 519948 105488 582820 105584
rect 1104 104944 68000 105040
rect 519948 104944 582820 105040
rect 1104 104400 68000 104496
rect 519948 104400 582820 104496
rect 1104 103856 68000 103952
rect 519948 103856 582820 103952
rect 1104 103312 68000 103408
rect 519948 103312 582820 103408
rect 1104 102768 68000 102864
rect 519948 102768 582820 102864
rect 1104 102224 68000 102320
rect 519948 102224 582820 102320
rect 1104 101680 68000 101776
rect 519948 101680 582820 101776
rect 1104 101136 68000 101232
rect 519948 101136 582820 101232
rect 1104 100592 68000 100688
rect 519948 100592 582820 100688
rect 520918 100512 520924 100564
rect 520976 100552 520982 100564
rect 580166 100552 580172 100564
rect 520976 100524 580172 100552
rect 520976 100512 520982 100524
rect 580166 100512 580172 100524
rect 580224 100512 580230 100564
rect 1104 100048 68000 100144
rect 519948 100048 582820 100144
rect 1104 99504 68000 99600
rect 519948 99504 582820 99600
rect 1104 98960 68000 99056
rect 519948 98960 582820 99056
rect 1104 98416 68000 98512
rect 519948 98416 582820 98512
rect 3510 97996 3516 98048
rect 3568 98036 3574 98048
rect 67174 98036 67180 98048
rect 3568 98008 67180 98036
rect 3568 97996 3574 98008
rect 67174 97996 67180 98008
rect 67232 97996 67238 98048
rect 1104 97872 68000 97968
rect 519948 97872 582820 97968
rect 1104 97328 68000 97424
rect 519948 97328 582820 97424
rect 1104 96784 68000 96880
rect 519948 96784 582820 96880
rect 1104 96240 68000 96336
rect 519948 96240 582820 96336
rect 1104 95696 68000 95792
rect 519948 95696 582820 95792
rect 1104 95152 68000 95248
rect 519948 95152 582820 95248
rect 1104 94608 68000 94704
rect 519948 94608 582820 94704
rect 1104 94064 68000 94160
rect 519948 94064 582820 94160
rect 1104 93520 68000 93616
rect 519948 93520 582820 93616
rect 1104 92976 68000 93072
rect 519948 92976 582820 93072
rect 1104 92432 68000 92528
rect 519948 92432 582820 92528
rect 1104 91888 68000 91984
rect 519948 91888 582820 91984
rect 1104 91344 68000 91440
rect 519948 91344 582820 91440
rect 1104 90800 68000 90896
rect 519948 90800 582820 90896
rect 1104 90256 68000 90352
rect 519948 90256 582820 90352
rect 1104 89712 68000 89808
rect 519948 89712 582820 89808
rect 1104 89168 68000 89264
rect 519948 89168 582820 89264
rect 1104 88624 68000 88720
rect 519948 88624 582820 88720
rect 3418 88340 3424 88392
rect 3476 88380 3482 88392
rect 67450 88380 67456 88392
rect 3476 88352 67456 88380
rect 3476 88340 3482 88352
rect 67450 88340 67456 88352
rect 67508 88340 67514 88392
rect 1104 88080 68000 88176
rect 519948 88080 582820 88176
rect 73154 87796 73160 87848
rect 73212 87836 73218 87848
rect 74430 87836 74436 87848
rect 73212 87808 74436 87836
rect 73212 87796 73218 87808
rect 74430 87796 74436 87808
rect 74488 87796 74494 87848
rect 78674 87796 78680 87848
rect 78732 87836 78738 87848
rect 79950 87836 79956 87848
rect 78732 87808 79956 87836
rect 78732 87796 78738 87808
rect 79950 87796 79956 87808
rect 80008 87796 80014 87848
rect 110414 87796 110420 87848
rect 110472 87836 110478 87848
rect 111690 87836 111696 87848
rect 110472 87808 111696 87836
rect 110472 87796 110478 87808
rect 111690 87796 111696 87808
rect 111748 87796 111754 87848
rect 116026 87796 116032 87848
rect 116084 87836 116090 87848
rect 117210 87836 117216 87848
rect 116084 87808 117216 87836
rect 116084 87796 116090 87808
rect 117210 87796 117216 87808
rect 117268 87796 117274 87848
rect 147766 87796 147772 87848
rect 147824 87836 147830 87848
rect 148950 87836 148956 87848
rect 147824 87808 148956 87836
rect 147824 87796 147830 87808
rect 148950 87796 148956 87808
rect 149008 87796 149014 87848
rect 150526 87796 150532 87848
rect 150584 87836 150590 87848
rect 151710 87836 151716 87848
rect 150584 87808 151716 87836
rect 150584 87796 150590 87808
rect 151710 87796 151716 87808
rect 151768 87796 151774 87848
rect 158714 87796 158720 87848
rect 158772 87836 158778 87848
rect 159898 87836 159904 87848
rect 158772 87808 159904 87836
rect 158772 87796 158778 87808
rect 159898 87796 159904 87808
rect 159956 87796 159962 87848
rect 166994 87796 167000 87848
rect 167052 87836 167058 87848
rect 168086 87836 168092 87848
rect 167052 87808 168092 87836
rect 167052 87796 167058 87808
rect 168086 87796 168092 87808
rect 168144 87796 168150 87848
rect 169754 87796 169760 87848
rect 169812 87836 169818 87848
rect 170754 87836 170760 87848
rect 169812 87808 170760 87836
rect 169812 87796 169818 87808
rect 170754 87796 170760 87808
rect 170812 87796 170818 87848
rect 296714 87796 296720 87848
rect 296772 87836 296778 87848
rect 297990 87836 297996 87848
rect 296772 87808 297996 87836
rect 296772 87796 296778 87808
rect 297990 87796 297996 87808
rect 298048 87796 298054 87848
rect 299474 87796 299480 87848
rect 299532 87836 299538 87848
rect 300750 87836 300756 87848
rect 299532 87808 300756 87836
rect 299532 87796 299538 87808
rect 300750 87796 300756 87808
rect 300808 87796 300814 87848
rect 316034 87796 316040 87848
rect 316092 87836 316098 87848
rect 317034 87836 317040 87848
rect 316092 87808 317040 87836
rect 316092 87796 316098 87808
rect 317034 87796 317040 87808
rect 317092 87796 317098 87848
rect 321554 87796 321560 87848
rect 321612 87836 321618 87848
rect 322554 87836 322560 87848
rect 321612 87808 322560 87836
rect 321612 87796 321618 87808
rect 322554 87796 322560 87808
rect 322612 87796 322618 87848
rect 333974 87796 333980 87848
rect 334032 87836 334038 87848
rect 335250 87836 335256 87848
rect 334032 87808 335256 87836
rect 334032 87796 334038 87808
rect 335250 87796 335256 87808
rect 335308 87796 335314 87848
rect 402974 87796 402980 87848
rect 403032 87836 403038 87848
rect 404250 87836 404256 87848
rect 403032 87808 404256 87836
rect 403032 87796 403038 87808
rect 404250 87796 404256 87808
rect 404308 87796 404314 87848
rect 405734 87796 405740 87848
rect 405792 87836 405798 87848
rect 407010 87836 407016 87848
rect 405792 87808 407016 87836
rect 405792 87796 405798 87808
rect 407010 87796 407016 87808
rect 407068 87796 407074 87848
rect 408494 87796 408500 87848
rect 408552 87836 408558 87848
rect 409770 87836 409776 87848
rect 408552 87808 409776 87836
rect 408552 87796 408558 87808
rect 409770 87796 409776 87808
rect 409828 87796 409834 87848
rect 422294 87796 422300 87848
rect 422352 87836 422358 87848
rect 423386 87836 423392 87848
rect 422352 87808 423392 87836
rect 422352 87796 422358 87808
rect 423386 87796 423392 87808
rect 423444 87796 423450 87848
rect 430574 87796 430580 87848
rect 430632 87836 430638 87848
rect 431574 87836 431580 87848
rect 430632 87808 431580 87836
rect 430632 87796 430638 87808
rect 431574 87796 431580 87808
rect 431632 87796 431638 87848
rect 443086 87796 443092 87848
rect 443144 87836 443150 87848
rect 444270 87836 444276 87848
rect 443144 87808 444276 87836
rect 443144 87796 443150 87808
rect 444270 87796 444276 87808
rect 444328 87796 444334 87848
rect 448514 87796 448520 87848
rect 448572 87836 448578 87848
rect 449698 87836 449704 87848
rect 448572 87808 449704 87836
rect 448572 87796 448578 87808
rect 449698 87796 449704 87808
rect 449756 87796 449762 87848
rect 454034 87796 454040 87848
rect 454092 87836 454098 87848
rect 455126 87836 455132 87848
rect 454092 87808 455132 87836
rect 454092 87796 454098 87808
rect 455126 87796 455132 87808
rect 455184 87796 455190 87848
rect 456794 87796 456800 87848
rect 456852 87836 456858 87848
rect 457886 87836 457892 87848
rect 456852 87808 457892 87836
rect 456852 87796 456858 87808
rect 457886 87796 457892 87808
rect 457944 87796 457950 87848
rect 459646 87796 459652 87848
rect 459704 87836 459710 87848
rect 460646 87836 460652 87848
rect 459704 87808 460652 87836
rect 459704 87796 459710 87808
rect 460646 87796 460652 87808
rect 460704 87796 460710 87848
rect 1104 87536 68000 87632
rect 519948 87536 582820 87632
rect 1104 86992 68000 87088
rect 519948 86992 582820 87088
rect 521470 86912 521476 86964
rect 521528 86952 521534 86964
rect 580166 86952 580172 86964
rect 521528 86924 580172 86952
rect 521528 86912 521534 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 1104 86448 68000 86544
rect 519948 86448 582820 86544
rect 76006 86096 76012 86148
rect 76064 86136 76070 86148
rect 77202 86136 77208 86148
rect 76064 86108 77208 86136
rect 76064 86096 76070 86108
rect 77202 86096 77208 86108
rect 77260 86096 77266 86148
rect 103514 86096 103520 86148
rect 103572 86136 103578 86148
rect 104434 86136 104440 86148
rect 103572 86108 104440 86136
rect 103572 86096 103578 86108
rect 104434 86096 104440 86108
rect 104492 86096 104498 86148
rect 106274 86096 106280 86148
rect 106332 86136 106338 86148
rect 107194 86136 107200 86148
rect 106332 86108 107200 86136
rect 106332 86096 106338 86108
rect 107194 86096 107200 86108
rect 107252 86096 107258 86148
rect 109034 86096 109040 86148
rect 109092 86136 109098 86148
rect 109954 86136 109960 86148
rect 109092 86108 109960 86136
rect 109092 86096 109098 86108
rect 109954 86096 109960 86108
rect 110012 86096 110018 86148
rect 140774 86096 140780 86148
rect 140832 86136 140838 86148
rect 141694 86136 141700 86148
rect 140832 86108 141700 86136
rect 140832 86096 140838 86108
rect 141694 86096 141700 86108
rect 141752 86096 141758 86148
rect 294046 86096 294052 86148
rect 294104 86136 294110 86148
rect 295242 86136 295248 86148
rect 294104 86108 295248 86136
rect 294104 86096 294110 86108
rect 295242 86096 295248 86108
rect 295300 86096 295306 86148
rect 331306 86096 331312 86148
rect 331364 86136 331370 86148
rect 332502 86136 332508 86148
rect 331364 86108 332508 86136
rect 331364 86096 331370 86108
rect 332502 86096 332508 86108
rect 332560 86096 332566 86148
rect 438854 86096 438860 86148
rect 438912 86136 438918 86148
rect 439774 86136 439780 86148
rect 438912 86108 439780 86136
rect 438912 86096 438918 86108
rect 439774 86096 439780 86108
rect 439832 86096 439838 86148
rect 445846 86096 445852 86148
rect 445904 86136 445910 86148
rect 447042 86136 447048 86148
rect 445904 86108 447048 86136
rect 445904 86096 445910 86108
rect 447042 86096 447048 86108
rect 447100 86096 447106 86148
rect 1104 85904 582820 86000
rect 76558 85484 76564 85536
rect 76616 85524 76622 85536
rect 78122 85524 78128 85536
rect 76616 85496 78128 85524
rect 76616 85484 76622 85496
rect 78122 85484 78128 85496
rect 78180 85484 78186 85536
rect 79318 85484 79324 85536
rect 79376 85524 79382 85536
rect 80882 85524 80888 85536
rect 79376 85496 80888 85524
rect 79376 85484 79382 85496
rect 80882 85484 80888 85496
rect 80940 85484 80946 85536
rect 94498 85484 94504 85536
rect 94556 85524 94562 85536
rect 95142 85524 95148 85536
rect 94556 85496 95148 85524
rect 94556 85484 94562 85496
rect 95142 85484 95148 85496
rect 95200 85484 95206 85536
rect 95418 85484 95424 85536
rect 95476 85524 95482 85536
rect 96430 85524 96436 85536
rect 95476 85496 96436 85524
rect 95476 85484 95482 85496
rect 96430 85484 96436 85496
rect 96488 85484 96494 85536
rect 97166 85484 97172 85536
rect 97224 85524 97230 85536
rect 97902 85524 97908 85536
rect 97224 85496 97908 85524
rect 97224 85484 97230 85496
rect 97902 85484 97908 85496
rect 97960 85484 97966 85536
rect 98086 85484 98092 85536
rect 98144 85524 98150 85536
rect 99282 85524 99288 85536
rect 98144 85496 99288 85524
rect 98144 85484 98150 85496
rect 99282 85484 99288 85496
rect 99340 85484 99346 85536
rect 99926 85484 99932 85536
rect 99984 85524 99990 85536
rect 100662 85524 100668 85536
rect 99984 85496 100668 85524
rect 99984 85484 99990 85496
rect 100662 85484 100668 85496
rect 100720 85484 100726 85536
rect 100846 85484 100852 85536
rect 100904 85524 100910 85536
rect 102042 85524 102048 85536
rect 100904 85496 102048 85524
rect 100904 85484 100910 85496
rect 102042 85484 102048 85496
rect 102100 85484 102106 85536
rect 115198 85484 115204 85536
rect 115256 85524 115262 85536
rect 116302 85524 116308 85536
rect 115256 85496 116308 85524
rect 115256 85484 115262 85496
rect 116302 85484 116308 85496
rect 116360 85484 116366 85536
rect 119338 85484 119344 85536
rect 119396 85524 119402 85536
rect 120810 85524 120816 85536
rect 119396 85496 120816 85524
rect 119396 85484 119402 85496
rect 120810 85484 120816 85496
rect 120868 85484 120874 85536
rect 130378 85484 130384 85536
rect 130436 85524 130442 85536
rect 131758 85524 131764 85536
rect 130436 85496 131764 85524
rect 130436 85484 130442 85496
rect 131758 85484 131764 85496
rect 131816 85484 131822 85536
rect 146938 85484 146944 85536
rect 146996 85524 147002 85536
rect 148042 85524 148048 85536
rect 146996 85496 148048 85524
rect 146996 85484 147002 85496
rect 148042 85484 148048 85496
rect 148100 85484 148106 85536
rect 176010 85484 176016 85536
rect 176068 85524 176074 85536
rect 177114 85524 177120 85536
rect 176068 85496 177120 85524
rect 176068 85484 176074 85496
rect 177114 85484 177120 85496
rect 177172 85484 177178 85536
rect 180794 85484 180800 85536
rect 180852 85524 180858 85536
rect 182174 85524 182180 85536
rect 180852 85496 182180 85524
rect 180852 85484 180858 85496
rect 182174 85484 182180 85496
rect 182232 85484 182238 85536
rect 182634 85484 182640 85536
rect 182692 85524 182698 85536
rect 184198 85524 184204 85536
rect 182692 85496 184204 85524
rect 182692 85484 182698 85496
rect 184198 85484 184204 85496
rect 184256 85484 184262 85536
rect 184382 85484 184388 85536
rect 184440 85524 184446 85536
rect 186958 85524 186964 85536
rect 184440 85496 186964 85524
rect 184440 85484 184446 85496
rect 186958 85484 186964 85496
rect 187016 85484 187022 85536
rect 187142 85484 187148 85536
rect 187200 85524 187206 85536
rect 187602 85524 187608 85536
rect 187200 85496 187608 85524
rect 187200 85484 187206 85496
rect 187602 85484 187608 85496
rect 187660 85484 187666 85536
rect 188062 85484 188068 85536
rect 188120 85524 188126 85536
rect 188982 85524 188988 85536
rect 188120 85496 188988 85524
rect 188120 85484 188126 85496
rect 188982 85484 188988 85496
rect 189040 85484 189046 85536
rect 190822 85484 190828 85536
rect 190880 85524 190886 85536
rect 191650 85524 191656 85536
rect 190880 85496 191656 85524
rect 190880 85484 190886 85496
rect 191650 85484 191656 85496
rect 191708 85484 191714 85536
rect 192570 85484 192576 85536
rect 192628 85524 192634 85536
rect 193122 85524 193128 85536
rect 192628 85496 193128 85524
rect 192628 85484 192634 85496
rect 193122 85484 193128 85496
rect 193180 85484 193186 85536
rect 193490 85484 193496 85536
rect 193548 85524 193554 85536
rect 194502 85524 194508 85536
rect 193548 85496 194508 85524
rect 193548 85484 193554 85496
rect 194502 85484 194508 85496
rect 194560 85484 194566 85536
rect 195330 85484 195336 85536
rect 195388 85524 195394 85536
rect 195882 85524 195888 85536
rect 195388 85496 195888 85524
rect 195388 85484 195394 85496
rect 195882 85484 195888 85496
rect 195940 85484 195946 85536
rect 196250 85484 196256 85536
rect 196308 85524 196314 85536
rect 197170 85524 197176 85536
rect 196308 85496 197176 85524
rect 196308 85484 196314 85496
rect 197170 85484 197176 85496
rect 197228 85484 197234 85536
rect 198090 85484 198096 85536
rect 198148 85524 198154 85536
rect 198642 85524 198648 85536
rect 198148 85496 198648 85524
rect 198148 85484 198154 85496
rect 198642 85484 198648 85496
rect 198700 85484 198706 85536
rect 198918 85484 198924 85536
rect 198976 85524 198982 85536
rect 199930 85524 199936 85536
rect 198976 85496 199936 85524
rect 198976 85484 198982 85496
rect 199930 85484 199936 85496
rect 199988 85484 199994 85536
rect 200758 85484 200764 85536
rect 200816 85524 200822 85536
rect 201402 85524 201408 85536
rect 200816 85496 201408 85524
rect 200816 85484 200822 85496
rect 201402 85484 201408 85496
rect 201460 85484 201466 85536
rect 201678 85484 201684 85536
rect 201736 85524 201742 85536
rect 202782 85524 202788 85536
rect 201736 85496 202788 85524
rect 201736 85484 201742 85496
rect 202782 85484 202788 85496
rect 202840 85484 202846 85536
rect 203518 85484 203524 85536
rect 203576 85524 203582 85536
rect 204162 85524 204168 85536
rect 203576 85496 204168 85524
rect 203576 85484 203582 85496
rect 204162 85484 204168 85496
rect 204220 85484 204226 85536
rect 204438 85484 204444 85536
rect 204496 85524 204502 85536
rect 205450 85524 205456 85536
rect 204496 85496 205456 85524
rect 204496 85484 204502 85496
rect 205450 85484 205456 85496
rect 205508 85484 205514 85536
rect 206186 85484 206192 85536
rect 206244 85524 206250 85536
rect 206922 85524 206928 85536
rect 206244 85496 206928 85524
rect 206244 85484 206250 85496
rect 206922 85484 206928 85496
rect 206980 85484 206986 85536
rect 208946 85484 208952 85536
rect 209004 85524 209010 85536
rect 209682 85524 209688 85536
rect 209004 85496 209688 85524
rect 209004 85484 209010 85496
rect 209682 85484 209688 85496
rect 209740 85484 209746 85536
rect 211706 85484 211712 85536
rect 211764 85524 211770 85536
rect 212442 85524 212448 85536
rect 211764 85496 212448 85524
rect 211764 85484 211770 85496
rect 212442 85484 212448 85496
rect 212500 85484 212506 85536
rect 212626 85484 212632 85536
rect 212684 85524 212690 85536
rect 213822 85524 213828 85536
rect 212684 85496 213828 85524
rect 212684 85484 212690 85496
rect 213822 85484 213828 85496
rect 213880 85484 213886 85536
rect 214374 85484 214380 85536
rect 214432 85524 214438 85536
rect 215202 85524 215208 85536
rect 214432 85496 215208 85524
rect 214432 85484 214438 85496
rect 215202 85484 215208 85496
rect 215260 85484 215266 85536
rect 215294 85484 215300 85536
rect 215352 85524 215358 85536
rect 216582 85524 216588 85536
rect 215352 85496 216588 85524
rect 215352 85484 215358 85496
rect 216582 85484 216588 85496
rect 216640 85484 216646 85536
rect 217134 85484 217140 85536
rect 217192 85524 217198 85536
rect 217962 85524 217968 85536
rect 217192 85496 217968 85524
rect 217192 85484 217198 85496
rect 217962 85484 217968 85496
rect 218020 85484 218026 85536
rect 218054 85484 218060 85536
rect 218112 85524 218118 85536
rect 219342 85524 219348 85536
rect 218112 85496 219348 85524
rect 218112 85484 218118 85496
rect 219342 85484 219348 85496
rect 219400 85484 219406 85536
rect 219894 85484 219900 85536
rect 219952 85524 219958 85536
rect 220722 85524 220728 85536
rect 219952 85496 220728 85524
rect 219952 85484 219958 85496
rect 220722 85484 220728 85496
rect 220780 85484 220786 85536
rect 222562 85484 222568 85536
rect 222620 85524 222626 85536
rect 223482 85524 223488 85536
rect 222620 85496 223488 85524
rect 222620 85484 222626 85496
rect 223482 85484 223488 85496
rect 223540 85484 223546 85536
rect 224402 85484 224408 85536
rect 224460 85524 224466 85536
rect 224862 85524 224868 85536
rect 224460 85496 224868 85524
rect 224460 85484 224466 85496
rect 224862 85484 224868 85496
rect 224920 85484 224926 85536
rect 225322 85484 225328 85536
rect 225380 85524 225386 85536
rect 226150 85524 226156 85536
rect 225380 85496 226156 85524
rect 225380 85484 225386 85496
rect 226150 85484 226156 85496
rect 226208 85484 226214 85536
rect 227162 85484 227168 85536
rect 227220 85524 227226 85536
rect 227622 85524 227628 85536
rect 227220 85496 227628 85524
rect 227220 85484 227226 85496
rect 227622 85484 227628 85496
rect 227680 85484 227686 85536
rect 229830 85484 229836 85536
rect 229888 85524 229894 85536
rect 230290 85524 230296 85536
rect 229888 85496 230296 85524
rect 229888 85484 229894 85496
rect 230290 85484 230296 85496
rect 230348 85484 230354 85536
rect 230750 85484 230756 85536
rect 230808 85524 230814 85536
rect 231762 85524 231768 85536
rect 230808 85496 231768 85524
rect 230808 85484 230814 85496
rect 231762 85484 231768 85496
rect 231820 85484 231826 85536
rect 232590 85484 232596 85536
rect 232648 85524 232654 85536
rect 233142 85524 233148 85536
rect 232648 85496 233148 85524
rect 232648 85484 232654 85496
rect 233142 85484 233148 85496
rect 233200 85484 233206 85536
rect 233510 85484 233516 85536
rect 233568 85524 233574 85536
rect 234430 85524 234436 85536
rect 233568 85496 234436 85524
rect 233568 85484 233574 85496
rect 234430 85484 234436 85496
rect 234488 85484 234494 85536
rect 235258 85484 235264 85536
rect 235316 85524 235322 85536
rect 235902 85524 235908 85536
rect 235316 85496 235908 85524
rect 235316 85484 235322 85496
rect 235902 85484 235908 85496
rect 235960 85484 235966 85536
rect 236178 85484 236184 85536
rect 236236 85524 236242 85536
rect 237190 85524 237196 85536
rect 236236 85496 237196 85524
rect 236236 85484 236242 85496
rect 237190 85484 237196 85496
rect 237248 85484 237254 85536
rect 238018 85484 238024 85536
rect 238076 85524 238082 85536
rect 238662 85524 238668 85536
rect 238076 85496 238668 85524
rect 238076 85484 238082 85496
rect 238662 85484 238668 85496
rect 238720 85484 238726 85536
rect 240778 85484 240784 85536
rect 240836 85524 240842 85536
rect 241330 85524 241336 85536
rect 240836 85496 241336 85524
rect 240836 85484 240842 85496
rect 241330 85484 241336 85496
rect 241388 85484 241394 85536
rect 241698 85484 241704 85536
rect 241756 85524 241762 85536
rect 242710 85524 242716 85536
rect 241756 85496 242716 85524
rect 241756 85484 241762 85496
rect 242710 85484 242716 85496
rect 242768 85484 242774 85536
rect 243446 85484 243452 85536
rect 243504 85524 243510 85536
rect 244182 85524 244188 85536
rect 243504 85496 244188 85524
rect 243504 85484 243510 85496
rect 244182 85484 244188 85496
rect 244240 85484 244246 85536
rect 244366 85484 244372 85536
rect 244424 85524 244430 85536
rect 245562 85524 245568 85536
rect 244424 85496 245568 85524
rect 244424 85484 244430 85496
rect 245562 85484 245568 85496
rect 245620 85484 245626 85536
rect 246206 85484 246212 85536
rect 246264 85524 246270 85536
rect 246942 85524 246948 85536
rect 246264 85496 246948 85524
rect 246264 85484 246270 85496
rect 246942 85484 246948 85496
rect 247000 85484 247006 85536
rect 247126 85484 247132 85536
rect 247184 85524 247190 85536
rect 248322 85524 248328 85536
rect 247184 85496 248328 85524
rect 247184 85484 247190 85496
rect 248322 85484 248328 85496
rect 248380 85484 248386 85536
rect 248966 85484 248972 85536
rect 249024 85524 249030 85536
rect 249702 85524 249708 85536
rect 249024 85496 249708 85524
rect 249024 85484 249030 85496
rect 249702 85484 249708 85496
rect 249760 85484 249766 85536
rect 249794 85484 249800 85536
rect 249852 85524 249858 85536
rect 251082 85524 251088 85536
rect 249852 85496 251088 85524
rect 249852 85484 249858 85496
rect 251082 85484 251088 85496
rect 251140 85484 251146 85536
rect 251634 85484 251640 85536
rect 251692 85524 251698 85536
rect 252462 85524 252468 85536
rect 251692 85496 252468 85524
rect 251692 85484 251698 85496
rect 252462 85484 252468 85496
rect 252520 85484 252526 85536
rect 252554 85484 252560 85536
rect 252612 85524 252618 85536
rect 253842 85524 253848 85536
rect 252612 85496 253848 85524
rect 252612 85484 252618 85496
rect 253842 85484 253848 85496
rect 253900 85484 253906 85536
rect 254394 85484 254400 85536
rect 254452 85524 254458 85536
rect 255222 85524 255228 85536
rect 254452 85496 255228 85524
rect 254452 85484 254458 85496
rect 255222 85484 255228 85496
rect 255280 85484 255286 85536
rect 255314 85484 255320 85536
rect 255372 85524 255378 85536
rect 256602 85524 256608 85536
rect 255372 85496 256608 85524
rect 255372 85484 255378 85496
rect 256602 85484 256608 85496
rect 256660 85484 256666 85536
rect 256694 85484 256700 85536
rect 256752 85524 256758 85536
rect 257982 85524 257988 85536
rect 256752 85496 257988 85524
rect 256752 85484 256758 85496
rect 257982 85484 257988 85496
rect 258040 85484 258046 85536
rect 258074 85484 258080 85536
rect 258132 85524 258138 85536
rect 258902 85524 258908 85536
rect 258132 85496 258908 85524
rect 258132 85484 258138 85496
rect 258902 85484 258908 85496
rect 258960 85484 258966 85536
rect 259822 85484 259828 85536
rect 259880 85524 259886 85536
rect 260742 85524 260748 85536
rect 259880 85496 260748 85524
rect 259880 85484 259886 85496
rect 260742 85484 260748 85496
rect 260800 85484 260806 85536
rect 262582 85484 262588 85536
rect 262640 85524 262646 85536
rect 263502 85524 263508 85536
rect 262640 85496 263508 85524
rect 262640 85484 262646 85496
rect 263502 85484 263508 85496
rect 263560 85484 263566 85536
rect 264330 85484 264336 85536
rect 264388 85524 264394 85536
rect 264882 85524 264888 85536
rect 264388 85496 264888 85524
rect 264388 85484 264394 85496
rect 264882 85484 264888 85496
rect 264940 85484 264946 85536
rect 265250 85484 265256 85536
rect 265308 85524 265314 85536
rect 266262 85524 266268 85536
rect 265308 85496 266268 85524
rect 265308 85484 265314 85496
rect 266262 85484 266268 85496
rect 266320 85484 266326 85536
rect 267090 85484 267096 85536
rect 267148 85524 267154 85536
rect 267642 85524 267648 85536
rect 267148 85496 267648 85524
rect 267148 85484 267154 85496
rect 267642 85484 267648 85496
rect 267700 85484 267706 85536
rect 268010 85484 268016 85536
rect 268068 85524 268074 85536
rect 269022 85524 269028 85536
rect 268068 85496 269028 85524
rect 268068 85484 268074 85496
rect 269022 85484 269028 85496
rect 269080 85484 269086 85536
rect 269850 85484 269856 85536
rect 269908 85524 269914 85536
rect 270402 85524 270408 85536
rect 269908 85496 270408 85524
rect 269908 85484 269914 85496
rect 270402 85484 270408 85496
rect 270460 85484 270466 85536
rect 270770 85484 270776 85536
rect 270828 85524 270834 85536
rect 271782 85524 271788 85536
rect 270828 85496 271788 85524
rect 270828 85484 270834 85496
rect 271782 85484 271788 85496
rect 271840 85484 271846 85536
rect 272518 85484 272524 85536
rect 272576 85524 272582 85536
rect 273162 85524 273168 85536
rect 272576 85496 273168 85524
rect 272576 85484 272582 85496
rect 273162 85484 273168 85496
rect 273220 85484 273226 85536
rect 273438 85484 273444 85536
rect 273496 85524 273502 85536
rect 274542 85524 274548 85536
rect 273496 85496 274548 85524
rect 273496 85484 273502 85496
rect 274542 85484 274548 85496
rect 274600 85484 274606 85536
rect 275278 85484 275284 85536
rect 275336 85524 275342 85536
rect 275922 85524 275928 85536
rect 275336 85496 275928 85524
rect 275336 85484 275342 85496
rect 275922 85484 275928 85496
rect 275980 85484 275986 85536
rect 276198 85484 276204 85536
rect 276256 85524 276262 85536
rect 277210 85524 277216 85536
rect 276256 85496 277216 85524
rect 276256 85484 276262 85496
rect 277210 85484 277216 85496
rect 277268 85484 277274 85536
rect 278038 85484 278044 85536
rect 278096 85524 278102 85536
rect 278682 85524 278688 85536
rect 278096 85496 278688 85524
rect 278096 85484 278102 85496
rect 278682 85484 278688 85496
rect 278740 85484 278746 85536
rect 278958 85484 278964 85536
rect 279016 85524 279022 85536
rect 280062 85524 280068 85536
rect 279016 85496 280068 85524
rect 279016 85484 279022 85496
rect 280062 85484 280068 85496
rect 280120 85484 280126 85536
rect 280154 85484 280160 85536
rect 280212 85524 280218 85536
rect 280706 85524 280712 85536
rect 280212 85496 280712 85524
rect 280212 85484 280218 85496
rect 280706 85484 280712 85496
rect 280764 85484 280770 85536
rect 280798 85484 280804 85536
rect 280856 85524 280862 85536
rect 282546 85524 282552 85536
rect 280856 85496 282552 85524
rect 280856 85484 280862 85496
rect 282546 85484 282552 85496
rect 282604 85484 282610 85536
rect 289078 85484 289084 85536
rect 289136 85524 289142 85536
rect 289814 85524 289820 85536
rect 289136 85496 289820 85524
rect 289136 85484 289142 85496
rect 289814 85484 289820 85496
rect 289872 85484 289878 85536
rect 308398 85484 308404 85536
rect 308456 85524 308462 85536
rect 309778 85524 309784 85536
rect 308456 85496 309784 85524
rect 308456 85484 308462 85496
rect 309778 85484 309784 85496
rect 309836 85484 309842 85536
rect 309870 85484 309876 85536
rect 309928 85524 309934 85536
rect 310698 85524 310704 85536
rect 309928 85496 310704 85524
rect 309928 85484 309934 85496
rect 310698 85484 310704 85496
rect 310756 85484 310762 85536
rect 312538 85484 312544 85536
rect 312596 85524 312602 85536
rect 313458 85524 313464 85536
rect 312596 85496 313464 85524
rect 312596 85484 312602 85496
rect 313458 85484 313464 85496
rect 313516 85484 313522 85536
rect 337102 85484 337108 85536
rect 337160 85524 337166 85536
rect 338022 85524 338028 85536
rect 337160 85496 338028 85524
rect 337160 85484 337166 85496
rect 338022 85484 338028 85496
rect 338080 85484 338086 85536
rect 338850 85484 338856 85536
rect 338908 85524 338914 85536
rect 339402 85524 339408 85536
rect 338908 85496 339408 85524
rect 338908 85484 338914 85496
rect 339402 85484 339408 85496
rect 339460 85484 339466 85536
rect 339770 85484 339776 85536
rect 339828 85524 339834 85536
rect 340782 85524 340788 85536
rect 339828 85496 340788 85524
rect 339828 85484 339834 85496
rect 340782 85484 340788 85496
rect 340840 85484 340846 85536
rect 341610 85484 341616 85536
rect 341668 85524 341674 85536
rect 342162 85524 342168 85536
rect 341668 85496 342168 85524
rect 341668 85484 341674 85496
rect 342162 85484 342168 85496
rect 342220 85484 342226 85536
rect 342530 85484 342536 85536
rect 342588 85524 342594 85536
rect 343450 85524 343456 85536
rect 342588 85496 343456 85524
rect 342588 85484 342594 85496
rect 343450 85484 343456 85496
rect 343508 85484 343514 85536
rect 344370 85484 344376 85536
rect 344428 85524 344434 85536
rect 344922 85524 344928 85536
rect 344428 85496 344928 85524
rect 344428 85484 344434 85496
rect 344922 85484 344928 85496
rect 344980 85484 344986 85536
rect 345198 85484 345204 85536
rect 345256 85524 345262 85536
rect 346302 85524 346308 85536
rect 345256 85496 346308 85524
rect 345256 85484 345262 85496
rect 346302 85484 346308 85496
rect 346360 85484 346366 85536
rect 347038 85484 347044 85536
rect 347096 85524 347102 85536
rect 347682 85524 347688 85536
rect 347096 85496 347688 85524
rect 347096 85484 347102 85496
rect 347682 85484 347688 85496
rect 347740 85484 347746 85536
rect 347958 85484 347964 85536
rect 348016 85524 348022 85536
rect 348970 85524 348976 85536
rect 348016 85496 348976 85524
rect 348016 85484 348022 85496
rect 348970 85484 348976 85496
rect 349028 85484 349034 85536
rect 349798 85484 349804 85536
rect 349856 85524 349862 85536
rect 350442 85524 350448 85536
rect 349856 85496 350448 85524
rect 349856 85484 349862 85496
rect 350442 85484 350448 85496
rect 350500 85484 350506 85536
rect 350718 85484 350724 85536
rect 350776 85524 350782 85536
rect 351822 85524 351828 85536
rect 350776 85496 351828 85524
rect 350776 85484 350782 85496
rect 351822 85484 351828 85496
rect 351880 85484 351886 85536
rect 353386 85484 353392 85536
rect 353444 85524 353450 85536
rect 354490 85524 354496 85536
rect 353444 85496 354496 85524
rect 353444 85484 353450 85496
rect 354490 85484 354496 85496
rect 354548 85484 354554 85536
rect 355226 85484 355232 85536
rect 355284 85524 355290 85536
rect 355962 85524 355968 85536
rect 355284 85496 355968 85524
rect 355284 85484 355290 85496
rect 355962 85484 355968 85496
rect 356020 85484 356026 85536
rect 356146 85484 356152 85536
rect 356204 85524 356210 85536
rect 357250 85524 357256 85536
rect 356204 85496 357256 85524
rect 356204 85484 356210 85496
rect 357250 85484 357256 85496
rect 357308 85484 357314 85536
rect 357986 85484 357992 85536
rect 358044 85524 358050 85536
rect 358722 85524 358728 85536
rect 358044 85496 358728 85524
rect 358044 85484 358050 85496
rect 358722 85484 358728 85496
rect 358780 85484 358786 85536
rect 358906 85484 358912 85536
rect 358964 85524 358970 85536
rect 360010 85524 360016 85536
rect 358964 85496 360016 85524
rect 358964 85484 358970 85496
rect 360010 85484 360016 85496
rect 360068 85484 360074 85536
rect 360654 85484 360660 85536
rect 360712 85524 360718 85536
rect 361482 85524 361488 85536
rect 360712 85496 361488 85524
rect 360712 85484 360718 85496
rect 361482 85484 361488 85496
rect 361540 85484 361546 85536
rect 361574 85484 361580 85536
rect 361632 85524 361638 85536
rect 362862 85524 362868 85536
rect 361632 85496 362868 85524
rect 361632 85484 361638 85496
rect 362862 85484 362868 85496
rect 362920 85484 362926 85536
rect 363414 85484 363420 85536
rect 363472 85524 363478 85536
rect 364242 85524 364248 85536
rect 363472 85496 364248 85524
rect 363472 85484 363478 85496
rect 364242 85484 364248 85496
rect 364300 85484 364306 85536
rect 364334 85484 364340 85536
rect 364392 85524 364398 85536
rect 365530 85524 365536 85536
rect 364392 85496 365536 85524
rect 364392 85484 364398 85496
rect 365530 85484 365536 85496
rect 365588 85484 365594 85536
rect 366174 85484 366180 85536
rect 366232 85524 366238 85536
rect 367002 85524 367008 85536
rect 366232 85496 367008 85524
rect 366232 85484 366238 85496
rect 367002 85484 367008 85496
rect 367060 85484 367066 85536
rect 367922 85484 367928 85536
rect 367980 85524 367986 85536
rect 368382 85524 368388 85536
rect 367980 85496 368388 85524
rect 367980 85484 367986 85496
rect 368382 85484 368388 85496
rect 368440 85484 368446 85536
rect 368842 85484 368848 85536
rect 368900 85524 368906 85536
rect 369762 85524 369768 85536
rect 368900 85496 369768 85524
rect 368900 85484 368906 85496
rect 369762 85484 369768 85496
rect 369820 85484 369826 85536
rect 370682 85484 370688 85536
rect 370740 85524 370746 85536
rect 371142 85524 371148 85536
rect 370740 85496 371148 85524
rect 370740 85484 370746 85496
rect 371142 85484 371148 85496
rect 371200 85484 371206 85536
rect 371602 85484 371608 85536
rect 371660 85524 371666 85536
rect 372430 85524 372436 85536
rect 371660 85496 372436 85524
rect 371660 85484 371666 85496
rect 372430 85484 372436 85496
rect 372488 85484 372494 85536
rect 374270 85484 374276 85536
rect 374328 85524 374334 85536
rect 375190 85524 375196 85536
rect 374328 85496 375196 85524
rect 374328 85484 374334 85496
rect 375190 85484 375196 85496
rect 375248 85484 375254 85536
rect 376110 85484 376116 85536
rect 376168 85524 376174 85536
rect 376662 85524 376668 85536
rect 376168 85496 376668 85524
rect 376168 85484 376174 85496
rect 376662 85484 376668 85496
rect 376720 85484 376726 85536
rect 377030 85484 377036 85536
rect 377088 85524 377094 85536
rect 378042 85524 378048 85536
rect 377088 85496 378048 85524
rect 377088 85484 377094 85496
rect 378042 85484 378048 85496
rect 378100 85484 378106 85536
rect 378870 85484 378876 85536
rect 378928 85524 378934 85536
rect 379422 85524 379428 85536
rect 378928 85496 379428 85524
rect 378928 85484 378934 85496
rect 379422 85484 379428 85496
rect 379480 85484 379486 85536
rect 379790 85484 379796 85536
rect 379848 85524 379854 85536
rect 380802 85524 380808 85536
rect 379848 85496 380808 85524
rect 379848 85484 379854 85496
rect 380802 85484 380808 85496
rect 380860 85484 380866 85536
rect 381630 85484 381636 85536
rect 381688 85524 381694 85536
rect 382182 85524 382188 85536
rect 381688 85496 382188 85524
rect 381688 85484 381694 85496
rect 382182 85484 382188 85496
rect 382240 85484 382246 85536
rect 382458 85484 382464 85536
rect 382516 85524 382522 85536
rect 383470 85524 383476 85536
rect 382516 85496 383476 85524
rect 382516 85484 382522 85496
rect 383470 85484 383476 85496
rect 383528 85484 383534 85536
rect 384298 85484 384304 85536
rect 384356 85524 384362 85536
rect 384942 85524 384948 85536
rect 384356 85496 384948 85524
rect 384356 85484 384362 85496
rect 384942 85484 384948 85496
rect 385000 85484 385006 85536
rect 385218 85484 385224 85536
rect 385276 85524 385282 85536
rect 386230 85524 386236 85536
rect 385276 85496 386236 85524
rect 385276 85484 385282 85496
rect 386230 85484 386236 85496
rect 386288 85484 386294 85536
rect 387058 85484 387064 85536
rect 387116 85524 387122 85536
rect 387702 85524 387708 85536
rect 387116 85496 387708 85524
rect 387116 85484 387122 85496
rect 387702 85484 387708 85496
rect 387760 85484 387766 85536
rect 387978 85484 387984 85536
rect 388036 85524 388042 85536
rect 389082 85524 389088 85536
rect 388036 85496 389088 85524
rect 388036 85484 388042 85496
rect 389082 85484 389088 85496
rect 389140 85484 389146 85536
rect 389726 85484 389732 85536
rect 389784 85524 389790 85536
rect 390462 85524 390468 85536
rect 389784 85496 390468 85524
rect 389784 85484 389790 85496
rect 390462 85484 390468 85496
rect 390520 85484 390526 85536
rect 390646 85484 390652 85536
rect 390704 85524 390710 85536
rect 391842 85524 391848 85536
rect 390704 85496 391848 85524
rect 390704 85484 390710 85496
rect 391842 85484 391848 85496
rect 391900 85484 391906 85536
rect 392486 85484 392492 85536
rect 392544 85524 392550 85536
rect 393222 85524 393228 85536
rect 392544 85496 393228 85524
rect 392544 85484 392550 85496
rect 393222 85484 393228 85496
rect 393280 85484 393286 85536
rect 393406 85484 393412 85536
rect 393464 85524 393470 85536
rect 394602 85524 394608 85536
rect 393464 85496 394608 85524
rect 393464 85484 393470 85496
rect 394602 85484 394608 85496
rect 394660 85484 394666 85536
rect 395246 85484 395252 85536
rect 395304 85524 395310 85536
rect 395982 85524 395988 85536
rect 395304 85496 395988 85524
rect 395304 85484 395310 85496
rect 395982 85484 395988 85496
rect 396040 85484 396046 85536
rect 396166 85484 396172 85536
rect 396224 85524 396230 85536
rect 397270 85524 397276 85536
rect 396224 85496 397276 85524
rect 396224 85484 396230 85496
rect 397270 85484 397276 85496
rect 397328 85484 397334 85536
rect 397914 85484 397920 85536
rect 397972 85524 397978 85536
rect 398742 85524 398748 85536
rect 397972 85496 398748 85524
rect 397972 85484 397978 85496
rect 398742 85484 398748 85496
rect 398800 85484 398806 85536
rect 401502 85484 401508 85536
rect 401560 85524 401566 85536
rect 402514 85524 402520 85536
rect 401560 85496 402520 85524
rect 401560 85484 401566 85496
rect 402514 85484 402520 85496
rect 402572 85484 402578 85536
rect 435358 85484 435364 85536
rect 435416 85524 435422 85536
rect 436094 85524 436100 85536
rect 435416 85496 436100 85524
rect 435416 85484 435422 85496
rect 436094 85484 436100 85496
rect 436152 85484 436158 85536
rect 439498 85484 439504 85536
rect 439556 85524 439562 85536
rect 441522 85524 441528 85536
rect 439556 85496 441528 85524
rect 439556 85484 439562 85496
rect 441522 85484 441528 85496
rect 441580 85484 441586 85536
rect 442258 85484 442264 85536
rect 442316 85524 442322 85536
rect 443362 85524 443368 85536
rect 442316 85496 443368 85524
rect 442316 85484 442322 85496
rect 443362 85484 443368 85496
rect 443420 85484 443426 85536
rect 462222 85484 462228 85536
rect 462280 85524 462286 85536
rect 484302 85524 484308 85536
rect 462280 85496 484308 85524
rect 462280 85484 462286 85496
rect 484302 85484 484308 85496
rect 484360 85484 484366 85536
rect 493318 85484 493324 85536
rect 493376 85524 493382 85536
rect 493962 85524 493968 85536
rect 493376 85496 493968 85524
rect 493376 85484 493382 85496
rect 493962 85484 493968 85496
rect 494020 85484 494026 85536
rect 494238 85484 494244 85536
rect 494296 85524 494302 85536
rect 495342 85524 495348 85536
rect 494296 85496 495348 85524
rect 494296 85484 494302 85496
rect 495342 85484 495348 85496
rect 495400 85484 495406 85536
rect 496078 85484 496084 85536
rect 496136 85524 496142 85536
rect 496722 85524 496728 85536
rect 496136 85496 496728 85524
rect 496136 85484 496142 85496
rect 496722 85484 496728 85496
rect 496780 85484 496786 85536
rect 496998 85484 497004 85536
rect 497056 85524 497062 85536
rect 498102 85524 498108 85536
rect 497056 85496 498108 85524
rect 497056 85484 497062 85496
rect 498102 85484 498108 85496
rect 498160 85484 498166 85536
rect 498838 85484 498844 85536
rect 498896 85524 498902 85536
rect 499482 85524 499488 85536
rect 498896 85496 499488 85524
rect 498896 85484 498902 85496
rect 499482 85484 499488 85496
rect 499540 85484 499546 85536
rect 499666 85484 499672 85536
rect 499724 85524 499730 85536
rect 500770 85524 500776 85536
rect 499724 85496 500776 85524
rect 499724 85484 499730 85496
rect 500770 85484 500776 85496
rect 500828 85484 500834 85536
rect 501506 85484 501512 85536
rect 501564 85524 501570 85536
rect 502242 85524 502248 85536
rect 501564 85496 502248 85524
rect 501564 85484 501570 85496
rect 502242 85484 502248 85496
rect 502300 85484 502306 85536
rect 502426 85484 502432 85536
rect 502484 85524 502490 85536
rect 503530 85524 503536 85536
rect 502484 85496 503536 85524
rect 502484 85484 502490 85496
rect 503530 85484 503536 85496
rect 503588 85484 503594 85536
rect 504266 85484 504272 85536
rect 504324 85524 504330 85536
rect 505002 85524 505008 85536
rect 504324 85496 505008 85524
rect 504324 85484 504330 85496
rect 505002 85484 505008 85496
rect 505060 85484 505066 85536
rect 505186 85484 505192 85536
rect 505244 85524 505250 85536
rect 506290 85524 506296 85536
rect 505244 85496 506296 85524
rect 505244 85484 505250 85496
rect 506290 85484 506296 85496
rect 506348 85484 506354 85536
rect 506934 85484 506940 85536
rect 506992 85524 506998 85536
rect 507762 85524 507768 85536
rect 506992 85496 507768 85524
rect 506992 85484 506998 85496
rect 507762 85484 507768 85496
rect 507820 85484 507826 85536
rect 507854 85484 507860 85536
rect 507912 85524 507918 85536
rect 509050 85524 509056 85536
rect 507912 85496 509056 85524
rect 507912 85484 507918 85496
rect 509050 85484 509056 85496
rect 509108 85484 509114 85536
rect 509694 85484 509700 85536
rect 509752 85524 509758 85536
rect 510522 85524 510528 85536
rect 509752 85496 510528 85524
rect 509752 85484 509758 85496
rect 510522 85484 510528 85496
rect 510580 85484 510586 85536
rect 510614 85484 510620 85536
rect 510672 85524 510678 85536
rect 511810 85524 511816 85536
rect 510672 85496 511816 85524
rect 510672 85484 510678 85496
rect 511810 85484 511816 85496
rect 511868 85484 511874 85536
rect 512454 85484 512460 85536
rect 512512 85524 512518 85536
rect 513282 85524 513288 85536
rect 512512 85496 513288 85524
rect 512512 85484 512518 85496
rect 513282 85484 513288 85496
rect 513340 85484 513346 85536
rect 514202 85484 514208 85536
rect 514260 85524 514266 85536
rect 514662 85524 514668 85536
rect 514260 85496 514668 85524
rect 514260 85484 514266 85496
rect 514662 85484 514668 85496
rect 514720 85484 514726 85536
rect 515122 85484 515128 85536
rect 515180 85524 515186 85536
rect 516042 85524 516048 85536
rect 515180 85496 516048 85524
rect 515180 85484 515186 85496
rect 516042 85484 516048 85496
rect 516100 85484 516106 85536
rect 516962 85484 516968 85536
rect 517020 85524 517026 85536
rect 517422 85524 517428 85536
rect 517020 85496 517428 85524
rect 517020 85484 517026 85496
rect 517422 85484 517428 85496
rect 517480 85484 517486 85536
rect 517882 85484 517888 85536
rect 517940 85524 517946 85536
rect 518802 85524 518808 85536
rect 517940 85496 518808 85524
rect 517940 85484 517946 85496
rect 518802 85484 518808 85496
rect 518860 85484 518866 85536
rect 1104 85360 582820 85456
rect 175918 85280 175924 85332
rect 175976 85320 175982 85332
rect 178034 85320 178040 85332
rect 175976 85292 178040 85320
rect 175976 85280 175982 85292
rect 178034 85280 178040 85292
rect 178092 85280 178098 85332
rect 183554 85280 183560 85332
rect 183612 85320 183618 85332
rect 184842 85320 184848 85332
rect 183612 85292 184848 85320
rect 183612 85280 183618 85292
rect 184842 85280 184848 85292
rect 184900 85280 184906 85332
rect 207106 85280 207112 85332
rect 207164 85320 207170 85332
rect 209038 85320 209044 85332
rect 207164 85292 209044 85320
rect 207164 85280 207170 85292
rect 209038 85280 209044 85292
rect 209096 85280 209102 85332
rect 209866 85280 209872 85332
rect 209924 85320 209930 85332
rect 214558 85320 214564 85332
rect 209924 85292 214564 85320
rect 209924 85280 209930 85292
rect 214558 85280 214564 85292
rect 214616 85280 214622 85332
rect 221642 85280 221648 85332
rect 221700 85320 221706 85332
rect 224218 85320 224224 85332
rect 221700 85292 224224 85320
rect 221700 85280 221706 85292
rect 224218 85280 224224 85292
rect 224276 85280 224282 85332
rect 238938 85280 238944 85332
rect 238996 85320 239002 85332
rect 240778 85320 240784 85332
rect 238996 85292 240784 85320
rect 238996 85280 239002 85292
rect 240778 85280 240784 85292
rect 240836 85280 240842 85332
rect 261662 85280 261668 85332
rect 261720 85320 261726 85332
rect 266998 85320 267004 85332
rect 261720 85292 267004 85320
rect 261720 85280 261726 85292
rect 266998 85280 267004 85292
rect 267056 85280 267062 85332
rect 279786 85280 279792 85332
rect 279844 85320 279850 85332
rect 280890 85320 280896 85332
rect 279844 85292 280896 85320
rect 279844 85280 279850 85292
rect 280890 85280 280896 85292
rect 280948 85280 280954 85332
rect 281626 85280 281632 85332
rect 281684 85320 281690 85332
rect 286410 85320 286416 85332
rect 281684 85292 286416 85320
rect 281684 85280 281690 85292
rect 286410 85280 286416 85292
rect 286468 85280 286474 85332
rect 310422 85280 310428 85332
rect 310480 85320 310486 85332
rect 311618 85320 311624 85332
rect 310480 85292 311624 85320
rect 310480 85280 310486 85292
rect 311618 85280 311624 85292
rect 311676 85280 311682 85332
rect 351638 85280 351644 85332
rect 351696 85320 351702 85332
rect 352650 85320 352656 85332
rect 351696 85292 352656 85320
rect 351696 85280 351702 85292
rect 352650 85280 352656 85292
rect 352708 85280 352714 85332
rect 455322 85280 455328 85332
rect 455380 85320 455386 85332
rect 482462 85320 482468 85332
rect 455380 85292 482468 85320
rect 455380 85280 455386 85292
rect 482462 85280 482468 85292
rect 482520 85280 482526 85332
rect 482922 85280 482928 85332
rect 482980 85320 482986 85332
rect 489730 85320 489736 85332
rect 482980 85292 489736 85320
rect 482980 85280 482986 85292
rect 489730 85280 489736 85292
rect 489788 85280 489794 85332
rect 513374 85280 513380 85332
rect 513432 85320 513438 85332
rect 514570 85320 514576 85332
rect 513432 85292 514576 85320
rect 513432 85280 513438 85292
rect 514570 85280 514576 85292
rect 514628 85280 514634 85332
rect 107562 85212 107568 85264
rect 107620 85252 107626 85264
rect 155310 85252 155316 85264
rect 107620 85224 155316 85252
rect 107620 85212 107626 85224
rect 155310 85212 155316 85224
rect 155368 85212 155374 85264
rect 451182 85212 451188 85264
rect 451240 85252 451246 85264
rect 481542 85252 481548 85264
rect 451240 85224 481548 85252
rect 451240 85212 451246 85224
rect 481542 85212 481548 85224
rect 481600 85212 481606 85264
rect 96522 85144 96528 85196
rect 96580 85184 96586 85196
rect 152642 85184 152648 85196
rect 96580 85156 152648 85184
rect 96580 85144 96586 85156
rect 152642 85144 152648 85156
rect 152700 85144 152706 85196
rect 161382 85144 161388 85196
rect 161440 85184 161446 85196
rect 175366 85184 175372 85196
rect 161440 85156 175372 85184
rect 161440 85144 161446 85156
rect 175366 85144 175372 85156
rect 175424 85144 175430 85196
rect 444282 85144 444288 85196
rect 444340 85184 444346 85196
rect 479702 85184 479708 85196
rect 444340 85156 479708 85184
rect 444340 85144 444346 85156
rect 479702 85144 479708 85156
rect 479760 85144 479766 85196
rect 18598 85076 18604 85128
rect 18656 85116 18662 85128
rect 132586 85116 132592 85128
rect 18656 85088 132592 85116
rect 18656 85076 18662 85088
rect 132586 85076 132592 85088
rect 132644 85076 132650 85128
rect 151722 85076 151728 85128
rect 151780 85116 151786 85128
rect 172606 85116 172612 85128
rect 151780 85088 172612 85116
rect 151780 85076 151786 85088
rect 172606 85076 172612 85088
rect 172664 85076 172670 85128
rect 437382 85076 437388 85128
rect 437440 85116 437446 85128
rect 477862 85116 477868 85128
rect 437440 85088 477868 85116
rect 437440 85076 437446 85088
rect 477862 85076 477868 85088
rect 477920 85076 477926 85128
rect 480162 85076 480168 85128
rect 480220 85116 480226 85128
rect 488810 85116 488816 85128
rect 480220 85088 488816 85116
rect 480220 85076 480226 85088
rect 488810 85076 488816 85088
rect 488868 85076 488874 85128
rect 19978 85008 19984 85060
rect 20036 85048 20042 85060
rect 161658 85048 161664 85060
rect 20036 85020 161664 85048
rect 20036 85008 20042 85020
rect 161658 85008 161664 85020
rect 161716 85008 161722 85060
rect 352466 85008 352472 85060
rect 352524 85048 352530 85060
rect 398098 85048 398104 85060
rect 352524 85020 398104 85048
rect 352524 85008 352530 85020
rect 398098 85008 398104 85020
rect 398156 85008 398162 85060
rect 423582 85008 423588 85060
rect 423640 85048 423646 85060
rect 474274 85048 474280 85060
rect 423640 85020 474280 85048
rect 423640 85008 423646 85020
rect 474274 85008 474280 85020
rect 474332 85008 474338 85060
rect 476022 85008 476028 85060
rect 476080 85048 476086 85060
rect 487890 85048 487896 85060
rect 476080 85020 487896 85048
rect 476080 85008 476086 85020
rect 487890 85008 487896 85020
rect 487948 85008 487954 85060
rect 7558 84940 7564 84992
rect 7616 84980 7622 84992
rect 165338 84980 165344 84992
rect 7616 84952 165344 84980
rect 7616 84940 7622 84952
rect 165338 84940 165344 84952
rect 165396 84940 165402 84992
rect 165522 84940 165528 84992
rect 165580 84980 165586 84992
rect 176286 84980 176292 84992
rect 165580 84952 176292 84980
rect 165580 84940 165586 84952
rect 176286 84940 176292 84952
rect 176344 84940 176350 84992
rect 189902 84940 189908 84992
rect 189960 84980 189966 84992
rect 195238 84980 195244 84992
rect 189960 84952 195244 84980
rect 189960 84940 189966 84952
rect 195238 84940 195244 84952
rect 195296 84940 195302 84992
rect 228910 84940 228916 84992
rect 228968 84980 228974 84992
rect 232498 84980 232504 84992
rect 228968 84952 232504 84980
rect 228968 84940 228974 84952
rect 232498 84940 232504 84952
rect 232556 84940 232562 84992
rect 239858 84940 239864 84992
rect 239916 84980 239922 84992
rect 249058 84980 249064 84992
rect 239916 84952 249064 84980
rect 239916 84940 239922 84952
rect 249058 84940 249064 84952
rect 249116 84940 249122 84992
rect 254578 84940 254584 84992
rect 254636 84980 254642 84992
rect 286226 84980 286232 84992
rect 254636 84952 286232 84980
rect 254636 84940 254642 84952
rect 286226 84940 286232 84952
rect 286284 84940 286290 84992
rect 287698 84940 287704 84992
rect 287756 84980 287762 84992
rect 401594 84980 401600 84992
rect 287756 84952 401600 84980
rect 287756 84940 287762 84952
rect 401594 84940 401600 84952
rect 401652 84940 401658 84992
rect 416682 84940 416688 84992
rect 416740 84980 416746 84992
rect 472434 84980 472440 84992
rect 416740 84952 472440 84980
rect 416740 84940 416746 84952
rect 472434 84940 472440 84952
rect 472492 84940 472498 84992
rect 473262 84940 473268 84992
rect 473320 84980 473326 84992
rect 486970 84980 486976 84992
rect 473320 84952 486976 84980
rect 473320 84940 473326 84952
rect 486970 84940 486976 84952
rect 487028 84940 487034 84992
rect 495158 84940 495164 84992
rect 495216 84980 495222 84992
rect 503806 84980 503812 84992
rect 495216 84952 503812 84980
rect 495216 84940 495222 84952
rect 503806 84940 503812 84952
rect 503864 84940 503870 84992
rect 1104 84816 582820 84912
rect 466362 84736 466368 84788
rect 466420 84776 466426 84788
rect 485130 84776 485136 84788
rect 466420 84748 485136 84776
rect 466420 84736 466426 84748
rect 485130 84736 485136 84748
rect 485188 84736 485194 84788
rect 469122 84668 469128 84720
rect 469180 84708 469186 84720
rect 486050 84708 486056 84720
rect 469180 84680 486056 84708
rect 469180 84668 469186 84680
rect 486050 84668 486056 84680
rect 486108 84668 486114 84720
rect 227990 84600 227996 84652
rect 228048 84640 228054 84652
rect 229738 84640 229744 84652
rect 228048 84612 229744 84640
rect 228048 84600 228054 84612
rect 229738 84600 229744 84612
rect 229796 84600 229802 84652
rect 373442 84600 373448 84652
rect 373500 84640 373506 84652
rect 376018 84640 376024 84652
rect 373500 84612 376024 84640
rect 373500 84600 373506 84612
rect 376018 84600 376024 84612
rect 376076 84600 376082 84652
rect 208026 84396 208032 84448
rect 208084 84436 208090 84448
rect 211798 84436 211804 84448
rect 208084 84408 211804 84436
rect 208084 84396 208090 84408
rect 211798 84396 211804 84408
rect 211856 84396 211862 84448
rect 1104 84272 582820 84368
rect 112438 84192 112444 84244
rect 112496 84232 112502 84244
rect 114462 84232 114468 84244
rect 112496 84204 114468 84232
rect 112496 84192 112502 84204
rect 114462 84192 114468 84204
rect 114520 84192 114526 84244
rect 169018 84192 169024 84244
rect 169076 84232 169082 84244
rect 171686 84232 171692 84244
rect 169076 84204 171692 84232
rect 169076 84192 169082 84204
rect 171686 84192 171692 84204
rect 171744 84192 171750 84244
rect 257062 84192 257068 84244
rect 257120 84232 257126 84244
rect 258718 84232 258724 84244
rect 257120 84204 258724 84232
rect 257120 84192 257126 84204
rect 258718 84192 258724 84204
rect 258776 84192 258782 84244
rect 286318 84192 286324 84244
rect 286376 84232 286382 84244
rect 287054 84232 287060 84244
rect 286376 84204 287060 84232
rect 286376 84192 286382 84204
rect 287054 84192 287060 84204
rect 287112 84192 287118 84244
rect 487062 84192 487068 84244
rect 487120 84232 487126 84244
rect 490650 84232 490656 84244
rect 487120 84204 490656 84232
rect 487120 84192 487126 84204
rect 490650 84192 490656 84204
rect 490708 84192 490714 84244
rect 1104 83728 582820 83824
rect 62022 83512 62028 83564
rect 62080 83552 62086 83564
rect 84286 83552 84292 83564
rect 62080 83524 84292 83552
rect 62080 83512 62086 83524
rect 84286 83512 84292 83524
rect 84344 83512 84350 83564
rect 153102 83512 153108 83564
rect 153160 83552 153166 83564
rect 288434 83552 288440 83564
rect 153160 83524 288440 83552
rect 153160 83512 153166 83524
rect 288434 83512 288440 83524
rect 288492 83512 288498 83564
rect 292482 83512 292488 83564
rect 292540 83552 292546 83564
rect 440326 83552 440332 83564
rect 292540 83524 440332 83552
rect 292540 83512 292546 83524
rect 440326 83512 440332 83524
rect 440384 83512 440390 83564
rect 10318 83444 10324 83496
rect 10376 83484 10382 83496
rect 71866 83484 71872 83496
rect 10376 83456 71872 83484
rect 10376 83444 10382 83456
rect 71866 83444 71872 83456
rect 71924 83444 71930 83496
rect 129642 83444 129648 83496
rect 129700 83484 129706 83496
rect 167086 83484 167092 83496
rect 129700 83456 167092 83484
rect 129700 83444 129706 83456
rect 167086 83444 167092 83456
rect 167144 83444 167150 83496
rect 184934 83444 184940 83496
rect 184992 83484 184998 83496
rect 200114 83484 200120 83496
rect 184992 83456 200120 83484
rect 184992 83444 184998 83456
rect 200114 83444 200120 83456
rect 200172 83444 200178 83496
rect 256694 83444 256700 83496
rect 256752 83484 256758 83496
rect 483106 83484 483112 83496
rect 256752 83456 483112 83484
rect 256752 83444 256758 83456
rect 483106 83444 483112 83456
rect 483164 83444 483170 83496
rect 1104 83184 582820 83280
rect 1104 82640 582820 82736
rect 309778 82220 309784 82272
rect 309836 82260 309842 82272
rect 444374 82260 444380 82272
rect 309836 82232 444380 82260
rect 309836 82220 309842 82232
rect 444374 82220 444380 82232
rect 444432 82220 444438 82272
rect 1104 82096 582820 82192
rect 1104 81552 582820 81648
rect 1104 81008 582820 81104
rect 241422 80792 241428 80844
rect 241480 80832 241486 80844
rect 310422 80832 310428 80844
rect 241480 80804 310428 80832
rect 241480 80792 241486 80804
rect 310422 80792 310428 80804
rect 310480 80792 310486 80844
rect 59262 80724 59268 80776
rect 59320 80764 59326 80776
rect 84102 80764 84108 80776
rect 59320 80736 84108 80764
rect 59320 80724 59326 80736
rect 84102 80724 84108 80736
rect 84160 80724 84166 80776
rect 133782 80724 133788 80776
rect 133840 80764 133846 80776
rect 166994 80764 167000 80776
rect 133840 80736 167000 80764
rect 133840 80724 133846 80736
rect 166994 80724 167000 80736
rect 167052 80724 167058 80776
rect 258074 80724 258080 80776
rect 258132 80764 258138 80776
rect 487154 80764 487160 80776
rect 258132 80736 487160 80764
rect 258132 80724 258138 80736
rect 487154 80724 487160 80736
rect 487212 80724 487218 80776
rect 14458 80656 14464 80708
rect 14516 80696 14522 80708
rect 102134 80696 102140 80708
rect 14516 80668 102140 80696
rect 14516 80656 14522 80668
rect 102134 80656 102140 80668
rect 102192 80656 102198 80708
rect 143442 80656 143448 80708
rect 143500 80696 143506 80708
rect 401502 80696 401508 80708
rect 143500 80668 401508 80696
rect 143500 80656 143506 80668
rect 401502 80656 401508 80668
rect 401560 80656 401566 80708
rect 1104 80464 582820 80560
rect 1104 79920 582820 80016
rect 1104 79376 582820 79472
rect 344830 79296 344836 79348
rect 344888 79336 344894 79348
rect 454126 79336 454132 79348
rect 344888 79308 454132 79336
rect 344888 79296 344894 79308
rect 454126 79296 454132 79308
rect 454184 79296 454190 79348
rect 1104 78832 582820 78928
rect 1104 78288 582820 78384
rect 230382 78072 230388 78124
rect 230440 78112 230446 78124
rect 307846 78112 307852 78124
rect 230440 78084 307852 78112
rect 230440 78072 230446 78084
rect 307846 78072 307852 78084
rect 307904 78072 307910 78124
rect 70210 78004 70216 78056
rect 70268 78044 70274 78056
rect 116026 78044 116032 78056
rect 70268 78016 116032 78044
rect 70268 78004 70274 78016
rect 116026 78004 116032 78016
rect 116084 78004 116090 78056
rect 137922 78004 137928 78056
rect 137980 78044 137986 78056
rect 284386 78044 284392 78056
rect 137980 78016 284392 78044
rect 137980 78004 137986 78016
rect 284386 78004 284392 78016
rect 284444 78004 284450 78056
rect 352558 78004 352564 78056
rect 352616 78044 352622 78056
rect 455414 78044 455420 78056
rect 352616 78016 455420 78044
rect 352616 78004 352622 78016
rect 455414 78004 455420 78016
rect 455472 78004 455478 78056
rect 12342 77936 12348 77988
rect 12400 77976 12406 77988
rect 73246 77976 73252 77988
rect 12400 77948 73252 77976
rect 12400 77936 12406 77948
rect 73246 77936 73252 77948
rect 73304 77936 73310 77988
rect 280154 77936 280160 77988
rect 280212 77976 280218 77988
rect 572714 77976 572720 77988
rect 280212 77948 572720 77976
rect 280212 77936 280218 77948
rect 572714 77936 572720 77948
rect 572772 77936 572778 77988
rect 1104 77744 582820 77840
rect 1104 77200 582820 77296
rect 1104 76656 582820 76752
rect 281442 76508 281448 76560
rect 281500 76548 281506 76560
rect 437474 76548 437480 76560
rect 281500 76520 437480 76548
rect 281500 76508 281506 76520
rect 437474 76508 437480 76520
rect 437532 76508 437538 76560
rect 1104 76112 582820 76208
rect 1104 75568 582820 75664
rect 227530 75284 227536 75336
rect 227588 75324 227594 75336
rect 307754 75324 307760 75336
rect 227588 75296 307760 75324
rect 227588 75284 227594 75296
rect 307754 75284 307760 75296
rect 307812 75284 307818 75336
rect 30282 75216 30288 75268
rect 30340 75256 30346 75268
rect 76006 75256 76012 75268
rect 30340 75228 76012 75256
rect 30340 75216 30346 75228
rect 76006 75216 76012 75228
rect 76064 75216 76070 75268
rect 155862 75216 155868 75268
rect 155920 75256 155926 75268
rect 289078 75256 289084 75268
rect 155920 75228 289084 75256
rect 155920 75216 155926 75228
rect 289078 75216 289084 75228
rect 289136 75216 289142 75268
rect 75822 75148 75828 75200
rect 75880 75188 75886 75200
rect 146386 75188 146392 75200
rect 75880 75160 146392 75188
rect 75880 75148 75886 75160
rect 146386 75148 146392 75160
rect 146444 75148 146450 75200
rect 280890 75148 280896 75200
rect 280948 75188 280954 75200
rect 568574 75188 568580 75200
rect 280948 75160 568580 75188
rect 280948 75148 280954 75160
rect 568574 75148 568580 75160
rect 568632 75148 568638 75200
rect 1104 75024 582820 75120
rect 1104 74480 582820 74576
rect 224218 74060 224224 74112
rect 224276 74100 224282 74112
rect 340874 74100 340880 74112
rect 224276 74072 340880 74100
rect 224276 74060 224282 74072
rect 340874 74060 340880 74072
rect 340932 74060 340938 74112
rect 1104 73936 582820 74032
rect 148962 73856 148968 73908
rect 149020 73896 149026 73908
rect 287146 73896 287152 73908
rect 149020 73868 287152 73896
rect 149020 73856 149026 73868
rect 287146 73856 287152 73868
rect 287204 73856 287210 73908
rect 375190 73856 375196 73908
rect 375248 73896 375254 73908
rect 484394 73896 484400 73908
rect 375248 73868 484400 73896
rect 375248 73856 375254 73868
rect 484394 73856 484400 73868
rect 484452 73856 484458 73908
rect 34422 73788 34428 73840
rect 34480 73828 34486 73840
rect 76558 73828 76564 73840
rect 34480 73800 76564 73828
rect 34480 73788 34486 73800
rect 76558 73788 76564 73800
rect 76616 73788 76622 73840
rect 92382 73788 92388 73840
rect 92440 73828 92446 73840
rect 121546 73828 121552 73840
rect 92440 73800 121552 73828
rect 92440 73788 92446 73800
rect 121546 73788 121552 73800
rect 121604 73788 121610 73840
rect 274358 73788 274364 73840
rect 274416 73828 274422 73840
rect 435358 73828 435364 73840
rect 274416 73800 435364 73828
rect 274416 73788 274422 73800
rect 435358 73788 435364 73800
rect 435416 73788 435422 73840
rect 1104 73392 582820 73488
rect 521378 73108 521384 73160
rect 521436 73148 521442 73160
rect 580166 73148 580172 73160
rect 521436 73120 580172 73148
rect 521436 73108 521442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 1104 72848 582820 72944
rect 1104 72304 582820 72400
rect 1104 71760 582820 71856
rect 1104 71216 582820 71312
rect 220630 71068 220636 71120
rect 220688 71108 220694 71120
rect 338114 71108 338120 71120
rect 220688 71080 338120 71108
rect 220688 71068 220694 71080
rect 338114 71068 338120 71080
rect 338172 71068 338178 71120
rect 37182 71000 37188 71052
rect 37240 71040 37246 71052
rect 78766 71040 78772 71052
rect 37240 71012 78772 71040
rect 37240 71000 37246 71012
rect 78766 71000 78772 71012
rect 78824 71000 78830 71052
rect 255222 71000 255228 71052
rect 255280 71040 255286 71052
rect 469306 71040 469312 71052
rect 255280 71012 469312 71040
rect 255280 71000 255286 71012
rect 469306 71000 469312 71012
rect 469364 71000 469370 71052
rect 1104 70672 582820 70768
rect 1104 70128 582820 70224
rect 1104 69584 582820 69680
rect 1104 69040 582820 69136
rect 1104 68496 582820 68592
rect 220722 68348 220728 68400
rect 220780 68388 220786 68400
rect 334158 68388 334164 68400
rect 220780 68360 334164 68388
rect 220780 68348 220786 68360
rect 334158 68348 334164 68360
rect 334216 68348 334222 68400
rect 15838 68280 15844 68332
rect 15896 68320 15902 68332
rect 103606 68320 103612 68332
rect 15896 68292 103612 68320
rect 15896 68280 15902 68292
rect 103606 68280 103612 68292
rect 103664 68280 103670 68332
rect 253750 68280 253756 68332
rect 253808 68320 253814 68332
rect 465258 68320 465264 68332
rect 253808 68292 465264 68320
rect 253808 68280 253814 68292
rect 465258 68280 465264 68292
rect 465316 68280 465322 68332
rect 1104 67952 582820 68048
rect 1104 67408 582820 67504
rect 252278 66988 252284 67040
rect 252336 67028 252342 67040
rect 430666 67028 430672 67040
rect 252336 67000 430672 67028
rect 252336 66988 252342 67000
rect 430666 66988 430672 67000
rect 430724 66988 430730 67040
rect 1104 66864 582820 66960
rect 1104 66320 582820 66416
rect 1104 65776 582820 65872
rect 219250 65560 219256 65612
rect 219308 65600 219314 65612
rect 331398 65600 331404 65612
rect 219308 65572 331404 65600
rect 219308 65560 219314 65572
rect 331398 65560 331404 65572
rect 331456 65560 331462 65612
rect 349798 65560 349804 65612
rect 349856 65600 349862 65612
rect 454034 65600 454040 65612
rect 349856 65572 454040 65600
rect 349856 65560 349862 65572
rect 454034 65560 454040 65572
rect 454092 65560 454098 65612
rect 28902 65492 28908 65544
rect 28960 65532 28966 65544
rect 106366 65532 106372 65544
rect 28960 65504 106372 65532
rect 28960 65492 28966 65504
rect 106366 65492 106372 65504
rect 106424 65492 106430 65544
rect 252462 65492 252468 65544
rect 252520 65532 252526 65544
rect 458266 65532 458272 65544
rect 252520 65504 458272 65532
rect 252520 65492 252526 65504
rect 458266 65492 458272 65504
rect 458324 65492 458330 65544
rect 1104 65232 582820 65328
rect 1104 64688 582820 64784
rect 358078 64268 358084 64320
rect 358136 64308 358142 64320
rect 456886 64308 456892 64320
rect 358136 64280 456892 64308
rect 358136 64268 358142 64280
rect 456886 64268 456892 64280
rect 456944 64268 456950 64320
rect 1104 64144 582820 64240
rect 1104 63600 582820 63696
rect 1104 63056 582820 63152
rect 219342 62908 219348 62960
rect 219400 62948 219406 62960
rect 327258 62948 327264 62960
rect 219400 62920 327264 62948
rect 219400 62908 219406 62920
rect 327258 62908 327264 62920
rect 327316 62908 327322 62960
rect 324222 62840 324228 62892
rect 324280 62880 324286 62892
rect 448606 62880 448612 62892
rect 324280 62852 448612 62880
rect 324280 62840 324286 62852
rect 448606 62840 448612 62852
rect 448664 62840 448670 62892
rect 32398 62772 32404 62824
rect 32456 62812 32462 62824
rect 106274 62812 106280 62824
rect 32456 62784 106280 62812
rect 32456 62772 32462 62784
rect 106274 62772 106280 62784
rect 106332 62772 106338 62824
rect 241330 62772 241336 62824
rect 241388 62812 241394 62824
rect 415486 62812 415492 62824
rect 241388 62784 415492 62812
rect 241388 62772 241394 62784
rect 415486 62772 415492 62784
rect 415544 62772 415550 62824
rect 1104 62512 582820 62608
rect 1104 61968 582820 62064
rect 1104 61424 582820 61520
rect 146202 61344 146208 61396
rect 146260 61384 146266 61396
rect 403066 61384 403072 61396
rect 146260 61356 403072 61384
rect 146260 61344 146266 61356
rect 403066 61344 403072 61356
rect 403124 61344 403130 61396
rect 1104 60880 582820 60976
rect 521286 60664 521292 60716
rect 521344 60704 521350 60716
rect 580166 60704 580172 60716
rect 521344 60676 580172 60704
rect 521344 60664 521350 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 1104 60336 582820 60432
rect 217962 60120 217968 60172
rect 218020 60160 218026 60172
rect 324498 60160 324504 60172
rect 218020 60132 324504 60160
rect 218020 60120 218026 60132
rect 324498 60120 324504 60132
rect 324556 60120 324562 60172
rect 318058 60052 318064 60104
rect 318116 60092 318122 60104
rect 445846 60092 445852 60104
rect 318116 60064 445852 60092
rect 318116 60052 318122 60064
rect 445846 60052 445852 60064
rect 445904 60052 445910 60104
rect 38562 59984 38568 60036
rect 38620 60024 38626 60036
rect 109126 60024 109132 60036
rect 38620 59996 109132 60024
rect 38620 59984 38626 59996
rect 109126 59984 109132 59996
rect 109184 59984 109190 60036
rect 249058 59984 249064 60036
rect 249116 60024 249122 60036
rect 412726 60024 412732 60036
rect 249116 59996 412732 60024
rect 249116 59984 249122 59996
rect 412726 59984 412732 59996
rect 412784 59984 412790 60036
rect 1104 59792 582820 59888
rect 1104 59248 582820 59344
rect 1104 58704 582820 58800
rect 278038 58624 278044 58676
rect 278096 58664 278102 58676
rect 436186 58664 436192 58676
rect 278096 58636 436192 58664
rect 278096 58624 278102 58636
rect 436186 58624 436192 58636
rect 436244 58624 436250 58676
rect 1104 58160 582820 58256
rect 1104 57616 582820 57712
rect 216490 57332 216496 57384
rect 216548 57372 216554 57384
rect 320266 57372 320272 57384
rect 216548 57344 320272 57372
rect 216548 57332 216554 57344
rect 320266 57332 320272 57344
rect 320324 57332 320330 57384
rect 308490 57264 308496 57316
rect 308548 57304 308554 57316
rect 443086 57304 443092 57316
rect 308548 57276 443092 57304
rect 308548 57264 308554 57276
rect 443086 57264 443092 57276
rect 443144 57264 443150 57316
rect 10962 57196 10968 57248
rect 11020 57236 11026 57248
rect 130378 57236 130384 57248
rect 11020 57208 130384 57236
rect 11020 57196 11026 57208
rect 130378 57196 130384 57208
rect 130436 57196 130442 57248
rect 238662 57196 238668 57248
rect 238720 57236 238726 57248
rect 405918 57236 405924 57248
rect 238720 57208 405924 57236
rect 238720 57196 238726 57208
rect 405918 57196 405924 57208
rect 405976 57196 405982 57248
rect 1104 57072 582820 57168
rect 1104 56528 582820 56624
rect 216582 56108 216588 56160
rect 216640 56148 216646 56160
rect 316218 56148 316224 56160
rect 216640 56120 316224 56148
rect 216640 56108 216646 56120
rect 316218 56108 316224 56120
rect 316276 56108 316282 56160
rect 1104 55984 582820 56080
rect 299382 55904 299388 55956
rect 299440 55944 299446 55956
rect 441614 55944 441620 55956
rect 299440 55916 441620 55944
rect 299440 55904 299446 55916
rect 441614 55904 441620 55916
rect 441672 55904 441678 55956
rect 50982 55836 50988 55888
rect 51040 55876 51046 55888
rect 140866 55876 140872 55888
rect 51040 55848 140872 55876
rect 51040 55836 51046 55848
rect 140866 55836 140872 55848
rect 140924 55836 140930 55888
rect 237190 55836 237196 55888
rect 237248 55876 237254 55888
rect 399018 55876 399024 55888
rect 237248 55848 399024 55876
rect 237248 55836 237254 55848
rect 399018 55836 399024 55848
rect 399076 55836 399082 55888
rect 1104 55440 582820 55536
rect 1104 54896 582820 54992
rect 235810 54476 235816 54528
rect 235868 54516 235874 54528
rect 425146 54516 425152 54528
rect 235868 54488 425152 54516
rect 235868 54476 235874 54488
rect 425146 54476 425152 54488
rect 425204 54476 425210 54528
rect 1104 54352 582820 54448
rect 1104 53808 582820 53904
rect 1104 53264 582820 53360
rect 215202 53184 215208 53236
rect 215260 53224 215266 53236
rect 313366 53224 313372 53236
rect 215260 53196 313372 53224
rect 215260 53184 215266 53196
rect 313366 53184 313372 53196
rect 313424 53184 313430 53236
rect 285582 53116 285588 53168
rect 285640 53156 285646 53168
rect 438946 53156 438952 53168
rect 285640 53128 438952 53156
rect 285640 53116 285646 53128
rect 438946 53116 438952 53128
rect 439004 53116 439010 53168
rect 57882 53048 57888 53100
rect 57940 53088 57946 53100
rect 142154 53088 142160 53100
rect 57940 53060 142160 53088
rect 57940 53048 57946 53060
rect 142154 53048 142160 53060
rect 142212 53048 142218 53100
rect 235902 53048 235908 53100
rect 235960 53088 235966 53100
rect 394694 53088 394700 53100
rect 235960 53060 394700 53088
rect 235960 53048 235966 53060
rect 394694 53048 394700 53060
rect 394752 53048 394758 53100
rect 1104 52720 582820 52816
rect 1104 52176 582820 52272
rect 267550 51756 267556 51808
rect 267608 51796 267614 51808
rect 433426 51796 433432 51808
rect 267608 51768 433432 51796
rect 267608 51756 267614 51768
rect 433426 51756 433432 51768
rect 433484 51756 433490 51808
rect 1104 51632 582820 51728
rect 1104 51088 582820 51184
rect 1104 50544 582820 50640
rect 213730 50396 213736 50448
rect 213788 50436 213794 50448
rect 309134 50436 309140 50448
rect 213788 50408 309140 50436
rect 213788 50396 213794 50408
rect 309134 50396 309140 50408
rect 309192 50396 309198 50448
rect 377950 50396 377956 50448
rect 378008 50436 378014 50448
rect 485038 50436 485044 50448
rect 378008 50408 485044 50436
rect 378008 50396 378014 50408
rect 485038 50396 485044 50408
rect 485096 50396 485102 50448
rect 64782 50328 64788 50380
rect 64840 50368 64846 50380
rect 143626 50368 143632 50380
rect 64840 50340 143632 50368
rect 64840 50328 64846 50340
rect 143626 50328 143632 50340
rect 143684 50328 143690 50380
rect 234430 50328 234436 50380
rect 234488 50368 234494 50380
rect 387794 50368 387800 50380
rect 234488 50340 387800 50368
rect 234488 50328 234494 50340
rect 387794 50328 387800 50340
rect 387852 50328 387858 50380
rect 1104 50000 582820 50096
rect 1104 49456 582820 49552
rect 263318 49036 263324 49088
rect 263376 49076 263382 49088
rect 433334 49076 433340 49088
rect 263376 49048 433340 49076
rect 263376 49036 263382 49048
rect 433334 49036 433340 49048
rect 433392 49036 433398 49088
rect 1104 48912 582820 49008
rect 1104 48368 582820 48464
rect 1104 47824 582820 47920
rect 213822 47608 213828 47660
rect 213880 47648 213886 47660
rect 306466 47648 306472 47660
rect 213880 47620 306472 47648
rect 213880 47608 213886 47620
rect 306466 47608 306472 47620
rect 306524 47608 306530 47660
rect 378042 47608 378048 47660
rect 378100 47648 378106 47660
rect 487798 47648 487804 47660
rect 378100 47620 487804 47648
rect 378100 47608 378106 47620
rect 487798 47608 487804 47620
rect 487856 47608 487862 47660
rect 61930 47540 61936 47592
rect 61988 47580 61994 47592
rect 143534 47580 143540 47592
rect 61988 47552 143540 47580
rect 61988 47540 61994 47552
rect 143534 47540 143540 47552
rect 143592 47540 143598 47592
rect 233142 47540 233148 47592
rect 233200 47580 233206 47592
rect 383654 47580 383660 47592
rect 233200 47552 383660 47580
rect 233200 47540 233206 47552
rect 383654 47540 383660 47552
rect 383712 47540 383718 47592
rect 1104 47280 582820 47376
rect 521194 46860 521200 46912
rect 521252 46900 521258 46912
rect 580166 46900 580172 46912
rect 521252 46872 580172 46900
rect 521252 46860 521258 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 1104 46736 582820 46832
rect 256418 46316 256424 46368
rect 256476 46356 256482 46368
rect 430574 46356 430580 46368
rect 256476 46328 430580 46356
rect 256476 46316 256482 46328
rect 430574 46316 430580 46328
rect 430632 46316 430638 46368
rect 1104 46192 582820 46288
rect 1104 45648 582820 45744
rect 1104 45104 582820 45200
rect 344278 44956 344284 45008
rect 344336 44996 344342 45008
rect 452654 44996 452660 45008
rect 344336 44968 452660 44996
rect 344336 44956 344342 44968
rect 452654 44956 452660 44968
rect 452712 44956 452718 45008
rect 212442 44888 212448 44940
rect 212500 44928 212506 44940
rect 302418 44928 302424 44940
rect 212500 44900 302424 44928
rect 212500 44888 212506 44900
rect 302418 44888 302424 44900
rect 302476 44888 302482 44940
rect 376662 44888 376668 44940
rect 376720 44928 376726 44940
rect 489178 44928 489184 44940
rect 376720 44900 489184 44928
rect 376720 44888 376726 44900
rect 489178 44888 489184 44900
rect 489236 44888 489242 44940
rect 68922 44820 68928 44872
rect 68980 44860 68986 44872
rect 144914 44860 144920 44872
rect 68980 44832 144920 44860
rect 68980 44820 68986 44832
rect 144914 44820 144920 44832
rect 144972 44820 144978 44872
rect 231670 44820 231676 44872
rect 231728 44860 231734 44872
rect 380894 44860 380900 44872
rect 231728 44832 380900 44860
rect 231728 44820 231734 44832
rect 380894 44820 380900 44832
rect 380952 44820 380958 44872
rect 1104 44560 582820 44656
rect 1104 44016 582820 44112
rect 1104 43472 582820 43568
rect 231670 43392 231676 43444
rect 231728 43432 231734 43444
rect 425054 43432 425060 43444
rect 231728 43404 425060 43432
rect 231728 43392 231734 43404
rect 425054 43392 425060 43404
rect 425112 43392 425118 43444
rect 1104 42928 582820 43024
rect 1104 42384 582820 42480
rect 338758 42168 338764 42220
rect 338816 42208 338822 42220
rect 451366 42208 451372 42220
rect 338816 42180 451372 42208
rect 338816 42168 338822 42180
rect 451366 42168 451372 42180
rect 451424 42168 451430 42220
rect 211062 42100 211068 42152
rect 211120 42140 211126 42152
rect 299658 42140 299664 42152
rect 211120 42112 299664 42140
rect 211120 42100 211126 42112
rect 299658 42100 299664 42112
rect 299716 42100 299722 42152
rect 375282 42100 375288 42152
rect 375340 42140 375346 42152
rect 488534 42140 488540 42152
rect 375340 42112 488540 42140
rect 375340 42100 375346 42112
rect 488534 42100 488540 42112
rect 488592 42100 488598 42152
rect 53742 42032 53748 42084
rect 53800 42072 53806 42084
rect 140774 42072 140780 42084
rect 53800 42044 140780 42072
rect 53800 42032 53806 42044
rect 140774 42032 140780 42044
rect 140832 42032 140838 42084
rect 231762 42032 231768 42084
rect 231820 42072 231826 42084
rect 376754 42072 376760 42084
rect 231820 42044 376760 42072
rect 231820 42032 231826 42044
rect 376754 42032 376760 42044
rect 376812 42032 376818 42084
rect 1104 41840 582820 41936
rect 1104 41296 582820 41392
rect 1104 40752 582820 40848
rect 249610 40672 249616 40724
rect 249668 40712 249674 40724
rect 429194 40712 429200 40724
rect 249668 40684 429200 40712
rect 249668 40672 249674 40684
rect 429194 40672 429200 40684
rect 429252 40672 429258 40724
rect 1104 40208 582820 40304
rect 1104 39664 582820 39760
rect 214558 39380 214564 39432
rect 214616 39420 214622 39432
rect 295426 39420 295432 39432
rect 214616 39392 295432 39420
rect 214616 39380 214622 39392
rect 295426 39380 295432 39392
rect 295484 39380 295490 39432
rect 335998 39380 336004 39432
rect 336056 39420 336062 39432
rect 451274 39420 451280 39432
rect 336056 39392 451280 39420
rect 336056 39380 336062 39392
rect 451274 39380 451280 39392
rect 451332 39380 451338 39432
rect 71682 39312 71688 39364
rect 71740 39352 71746 39364
rect 146294 39352 146300 39364
rect 71740 39324 146300 39352
rect 71740 39312 71746 39324
rect 146294 39312 146300 39324
rect 146352 39312 146358 39364
rect 230290 39312 230296 39364
rect 230348 39352 230354 39364
rect 373994 39352 374000 39364
rect 230348 39324 374000 39352
rect 230348 39312 230354 39324
rect 373994 39312 374000 39324
rect 374052 39312 374058 39364
rect 376018 39312 376024 39364
rect 376076 39352 376082 39364
rect 481634 39352 481640 39364
rect 376076 39324 481640 39352
rect 376076 39312 376082 39324
rect 481634 39312 481640 39324
rect 481692 39312 481698 39364
rect 1104 39120 582820 39216
rect 1104 38576 582820 38672
rect 211798 38156 211804 38208
rect 211856 38196 211862 38208
rect 288434 38196 288440 38208
rect 211856 38168 288440 38196
rect 211856 38156 211862 38168
rect 288434 38156 288440 38168
rect 288492 38156 288498 38208
rect 1104 38032 582820 38128
rect 232498 37952 232504 38004
rect 232556 37992 232562 38004
rect 369854 37992 369860 38004
rect 232556 37964 369860 37992
rect 232556 37952 232562 37964
rect 369854 37952 369860 37964
rect 369912 37952 369918 38004
rect 35802 37884 35808 37936
rect 35860 37924 35866 37936
rect 107654 37924 107660 37936
rect 35860 37896 107660 37924
rect 35860 37884 35866 37896
rect 107654 37884 107660 37896
rect 107712 37884 107718 37936
rect 256510 37884 256516 37936
rect 256568 37924 256574 37936
rect 476298 37924 476304 37936
rect 256568 37896 476304 37924
rect 256568 37884 256574 37896
rect 476298 37884 476304 37896
rect 476356 37884 476362 37936
rect 1104 37488 582820 37584
rect 1104 36944 582820 37040
rect 245378 36524 245384 36576
rect 245436 36564 245442 36576
rect 427906 36564 427912 36576
rect 245436 36536 427912 36564
rect 245436 36524 245442 36536
rect 427906 36524 427912 36536
rect 427964 36524 427970 36576
rect 1104 36400 582820 36496
rect 1104 35856 582820 35952
rect 209038 35436 209044 35488
rect 209096 35476 209102 35488
rect 284478 35476 284484 35488
rect 209096 35448 284484 35476
rect 209096 35436 209102 35448
rect 284478 35436 284484 35448
rect 284536 35436 284542 35488
rect 1104 35312 582820 35408
rect 288342 35232 288348 35284
rect 288400 35272 288406 35284
rect 438854 35272 438860 35284
rect 288400 35244 438860 35272
rect 288400 35232 288406 35244
rect 438854 35232 438860 35244
rect 438912 35232 438918 35284
rect 45462 35164 45468 35216
rect 45520 35204 45526 35216
rect 110506 35204 110512 35216
rect 45520 35176 110512 35204
rect 45520 35164 45526 35176
rect 110506 35164 110512 35176
rect 110564 35164 110570 35216
rect 135162 35164 135168 35216
rect 135220 35204 135226 35216
rect 284294 35204 284300 35216
rect 135220 35176 284300 35204
rect 135220 35164 135226 35176
rect 284294 35164 284300 35176
rect 284352 35164 284358 35216
rect 286410 35164 286416 35216
rect 286468 35204 286474 35216
rect 575474 35204 575480 35216
rect 286468 35176 575480 35204
rect 286468 35164 286474 35176
rect 575474 35164 575480 35176
rect 575532 35164 575538 35216
rect 1104 34768 582820 34864
rect 1104 34224 582820 34320
rect 242618 33804 242624 33856
rect 242676 33844 242682 33856
rect 427814 33844 427820 33856
rect 242676 33816 427820 33844
rect 242676 33804 242682 33816
rect 427814 33804 427820 33816
rect 427872 33804 427878 33856
rect 1104 33680 582820 33776
rect 1104 33136 582820 33232
rect 521102 33056 521108 33108
rect 521160 33096 521166 33108
rect 580166 33096 580172 33108
rect 521160 33068 580172 33096
rect 521160 33056 521166 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 1104 32592 582820 32688
rect 206922 32512 206928 32564
rect 206980 32552 206986 32564
rect 281534 32552 281540 32564
rect 206980 32524 281540 32552
rect 206980 32512 206986 32524
rect 281534 32512 281540 32524
rect 281592 32512 281598 32564
rect 229738 32444 229744 32496
rect 229796 32484 229802 32496
rect 365714 32484 365720 32496
rect 229796 32456 365720 32484
rect 229796 32444 229802 32456
rect 365714 32444 365720 32456
rect 365772 32444 365778 32496
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 104894 32416 104900 32428
rect 23440 32388 104900 32416
rect 23440 32376 23446 32388
rect 104894 32376 104900 32388
rect 104952 32376 104958 32428
rect 117222 32376 117228 32428
rect 117280 32416 117286 32428
rect 128354 32416 128360 32428
rect 117280 32388 128360 32416
rect 117280 32376 117286 32388
rect 128354 32376 128360 32388
rect 128412 32376 128418 32428
rect 256602 32376 256608 32428
rect 256660 32416 256666 32428
rect 473446 32416 473452 32428
rect 256660 32388 473452 32416
rect 256660 32376 256666 32388
rect 473446 32376 473452 32388
rect 473504 32376 473510 32428
rect 1104 32048 582820 32144
rect 1104 31504 582820 31600
rect 237190 31084 237196 31136
rect 237248 31124 237254 31136
rect 309870 31124 309876 31136
rect 237248 31096 309876 31124
rect 237248 31084 237254 31096
rect 309870 31084 309876 31096
rect 309928 31084 309934 31136
rect 331122 31084 331128 31136
rect 331180 31124 331186 31136
rect 449894 31124 449900 31136
rect 331180 31096 449900 31124
rect 331180 31084 331186 31096
rect 449894 31084 449900 31096
rect 449952 31084 449958 31136
rect 1104 30960 582820 31056
rect 1104 30416 582820 30512
rect 1104 29872 582820 29968
rect 223298 29724 223304 29776
rect 223356 29764 223362 29776
rect 306374 29764 306380 29776
rect 223356 29736 306380 29764
rect 223356 29724 223362 29736
rect 306374 29724 306380 29736
rect 306432 29724 306438 29776
rect 144822 29656 144828 29708
rect 144880 29696 144886 29708
rect 286318 29696 286324 29708
rect 144880 29668 286324 29696
rect 144880 29656 144886 29668
rect 286318 29656 286324 29668
rect 286376 29656 286382 29708
rect 326982 29656 326988 29708
rect 327040 29696 327046 29708
rect 448514 29696 448520 29708
rect 327040 29668 448520 29696
rect 327040 29656 327046 29668
rect 448514 29656 448520 29668
rect 448572 29656 448578 29708
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 103514 29628 103520 29640
rect 19300 29600 103520 29628
rect 19300 29588 19306 29600
rect 103514 29588 103520 29600
rect 103572 29588 103578 29640
rect 113082 29588 113088 29640
rect 113140 29628 113146 29640
rect 127066 29628 127072 29640
rect 113140 29600 127072 29628
rect 113140 29588 113146 29600
rect 127066 29588 127072 29600
rect 127124 29588 127130 29640
rect 264882 29588 264888 29640
rect 264940 29628 264946 29640
rect 507854 29628 507860 29640
rect 264940 29600 507860 29628
rect 264940 29588 264946 29600
rect 507854 29588 507860 29600
rect 507912 29588 507918 29640
rect 1104 29328 582820 29424
rect 1104 28784 582820 28880
rect 248138 28364 248144 28416
rect 248196 28404 248202 28416
rect 312538 28404 312544 28416
rect 248196 28376 312544 28404
rect 248196 28364 248202 28376
rect 312538 28364 312544 28376
rect 312596 28364 312602 28416
rect 320818 28364 320824 28416
rect 320876 28404 320882 28416
rect 447134 28404 447140 28416
rect 320876 28376 447140 28404
rect 320876 28364 320882 28376
rect 447134 28364 447140 28376
rect 447192 28364 447198 28416
rect 1104 28240 582820 28336
rect 1104 27696 582820 27792
rect 1104 27152 582820 27248
rect 95050 26936 95056 26988
rect 95108 26976 95114 26988
rect 122834 26976 122840 26988
rect 95108 26948 122840 26976
rect 95108 26936 95114 26948
rect 122834 26936 122840 26948
rect 122892 26936 122898 26988
rect 162762 26936 162768 26988
rect 162820 26976 162826 26988
rect 291194 26976 291200 26988
rect 162820 26948 291200 26976
rect 162820 26936 162826 26948
rect 291194 26936 291200 26948
rect 291252 26936 291258 26988
rect 295242 26936 295248 26988
rect 295300 26976 295306 26988
rect 439498 26976 439504 26988
rect 295300 26948 439504 26976
rect 295300 26936 295306 26948
rect 439498 26936 439504 26948
rect 439556 26936 439562 26988
rect 42702 26868 42708 26920
rect 42760 26908 42766 26920
rect 109034 26908 109040 26920
rect 42760 26880 109040 26908
rect 42760 26868 42766 26880
rect 109034 26868 109040 26880
rect 109092 26868 109098 26920
rect 263410 26868 263416 26920
rect 263468 26908 263474 26920
rect 505094 26908 505100 26920
rect 263468 26880 505100 26908
rect 263468 26868 263474 26880
rect 505094 26868 505100 26880
rect 505152 26868 505158 26920
rect 1104 26608 582820 26704
rect 124122 26460 124128 26512
rect 124180 26500 124186 26512
rect 129826 26500 129832 26512
rect 124180 26472 129832 26500
rect 124180 26460 124186 26472
rect 129826 26460 129832 26472
rect 129884 26460 129890 26512
rect 1104 26064 582820 26160
rect 244090 25644 244096 25696
rect 244148 25684 244154 25696
rect 311894 25684 311900 25696
rect 244148 25656 311900 25684
rect 244148 25644 244154 25656
rect 311894 25644 311900 25656
rect 311952 25644 311958 25696
rect 313182 25644 313188 25696
rect 313240 25684 313246 25696
rect 445754 25684 445760 25696
rect 313240 25656 445760 25684
rect 313240 25644 313246 25656
rect 445754 25644 445760 25656
rect 445812 25644 445818 25696
rect 1104 25520 582820 25616
rect 1104 24976 582820 25072
rect 1104 24432 582820 24528
rect 128262 24216 128268 24268
rect 128320 24256 128326 24268
rect 280798 24256 280804 24268
rect 128320 24228 280804 24256
rect 128320 24216 128326 24228
rect 280798 24216 280804 24228
rect 280856 24216 280862 24268
rect 260558 24148 260564 24200
rect 260616 24188 260622 24200
rect 431954 24188 431960 24200
rect 260616 24160 431960 24188
rect 260616 24148 260622 24160
rect 431954 24148 431960 24160
rect 432012 24148 432018 24200
rect 88242 24080 88248 24132
rect 88300 24120 88306 24132
rect 121454 24120 121460 24132
rect 88300 24092 121460 24120
rect 88300 24080 88306 24092
rect 121454 24080 121460 24092
rect 121512 24080 121518 24132
rect 263502 24080 263508 24132
rect 263560 24120 263566 24132
rect 500954 24120 500960 24132
rect 263560 24092 500960 24120
rect 263560 24080 263566 24092
rect 500954 24080 500960 24092
rect 501012 24080 501018 24132
rect 1104 23888 582820 23984
rect 1104 23344 582820 23440
rect 234430 22924 234436 22976
rect 234488 22964 234494 22976
rect 308398 22964 308404 22976
rect 234488 22936 308404 22964
rect 234488 22924 234494 22936
rect 308398 22924 308404 22936
rect 308456 22924 308462 22976
rect 1104 22800 582820 22896
rect 302142 22720 302148 22772
rect 302200 22760 302206 22772
rect 442258 22760 442264 22772
rect 302200 22732 442264 22760
rect 302200 22720 302206 22732
rect 442258 22720 442264 22732
rect 442316 22720 442322 22772
rect 1104 22256 582820 22352
rect 1104 21712 582820 21808
rect 110322 21428 110328 21480
rect 110380 21468 110386 21480
rect 126974 21468 126980 21480
rect 110380 21440 126980 21468
rect 110380 21428 110386 21440
rect 126974 21428 126980 21440
rect 127032 21428 127038 21480
rect 147582 21428 147588 21480
rect 147640 21468 147646 21480
rect 169018 21468 169024 21480
rect 147640 21440 169024 21468
rect 147640 21428 147646 21440
rect 169018 21428 169024 21440
rect 169076 21428 169082 21480
rect 242710 21428 242716 21480
rect 242768 21468 242774 21480
rect 419718 21468 419724 21480
rect 242768 21440 419724 21468
rect 242768 21428 242774 21440
rect 419718 21428 419724 21440
rect 419776 21428 419782 21480
rect 53650 21360 53656 21412
rect 53708 21400 53714 21412
rect 111794 21400 111800 21412
rect 53708 21372 111800 21400
rect 53708 21360 53714 21372
rect 111794 21360 111800 21372
rect 111852 21360 111858 21412
rect 142062 21360 142068 21412
rect 142120 21400 142126 21412
rect 254578 21400 254584 21412
rect 142120 21372 254584 21400
rect 142120 21360 142126 21372
rect 254578 21360 254584 21372
rect 254636 21360 254642 21412
rect 266998 21360 267004 21412
rect 267056 21400 267062 21412
rect 498286 21400 498292 21412
rect 267056 21372 498292 21400
rect 267056 21360 267062 21372
rect 498286 21360 498292 21372
rect 498344 21360 498350 21412
rect 1104 21168 582820 21264
rect 1104 20624 582820 20720
rect 521010 20544 521016 20596
rect 521068 20584 521074 20596
rect 580166 20584 580172 20596
rect 521068 20556 580172 20584
rect 521068 20544 521074 20556
rect 580166 20544 580172 20556
rect 580224 20544 580230 20596
rect 1104 20080 582820 20176
rect 253842 19932 253848 19984
rect 253900 19972 253906 19984
rect 462498 19972 462504 19984
rect 253900 19944 462504 19972
rect 253900 19932 253906 19944
rect 462498 19932 462504 19944
rect 462556 19932 462562 19984
rect 1104 19536 582820 19632
rect 1104 18992 582820 19088
rect 160002 18708 160008 18760
rect 160060 18748 160066 18760
rect 289906 18748 289912 18760
rect 160060 18720 289912 18748
rect 160060 18708 160066 18720
rect 289906 18708 289912 18720
rect 289964 18708 289970 18760
rect 81342 18640 81348 18692
rect 81400 18680 81406 18692
rect 118786 18680 118792 18692
rect 81400 18652 118792 18680
rect 81400 18640 81406 18652
rect 118786 18640 118792 18652
rect 118844 18640 118850 18692
rect 140682 18640 140688 18692
rect 140740 18680 140746 18692
rect 169846 18680 169852 18692
rect 140740 18652 169852 18680
rect 140740 18640 140746 18652
rect 169846 18640 169852 18652
rect 169904 18640 169910 18692
rect 237282 18640 237288 18692
rect 237340 18680 237346 18692
rect 401594 18680 401600 18692
rect 237340 18652 401600 18680
rect 237340 18640 237346 18652
rect 401594 18640 401600 18652
rect 401652 18640 401658 18692
rect 45370 18572 45376 18624
rect 45428 18612 45434 18624
rect 79318 18612 79324 18624
rect 45428 18584 79324 18612
rect 45428 18572 45434 18584
rect 79318 18572 79324 18584
rect 79376 18572 79382 18624
rect 82722 18572 82728 18624
rect 82780 18612 82786 18624
rect 147766 18612 147772 18624
rect 82780 18584 147772 18612
rect 82780 18572 82786 18584
rect 147766 18572 147772 18584
rect 147824 18572 147830 18624
rect 188890 18572 188896 18624
rect 188948 18612 188954 18624
rect 213914 18612 213920 18624
rect 188948 18584 213920 18612
rect 188948 18572 188954 18584
rect 213914 18572 213920 18584
rect 213972 18572 213978 18624
rect 260650 18572 260656 18624
rect 260708 18612 260714 18624
rect 494054 18612 494060 18624
rect 260708 18584 494060 18612
rect 260708 18572 260714 18584
rect 494054 18572 494060 18584
rect 494112 18572 494118 18624
rect 1104 18448 582820 18544
rect 1104 17904 582820 18000
rect 1104 17360 582820 17456
rect 74442 17280 74448 17332
rect 74500 17320 74506 17332
rect 117314 17320 117320 17332
rect 74500 17292 117320 17320
rect 74500 17280 74506 17292
rect 117314 17280 117320 17292
rect 117372 17280 117378 17332
rect 144730 17280 144736 17332
rect 144788 17320 144794 17332
rect 169754 17320 169760 17332
rect 144788 17292 169760 17320
rect 144788 17280 144794 17292
rect 169754 17280 169760 17292
rect 169812 17280 169818 17332
rect 209682 17280 209688 17332
rect 209740 17320 209746 17332
rect 292758 17320 292764 17332
rect 209740 17292 292764 17320
rect 209740 17280 209746 17292
rect 292758 17280 292764 17292
rect 292816 17280 292822 17332
rect 352650 17280 352656 17332
rect 352708 17320 352714 17332
rect 396074 17320 396080 17332
rect 352708 17292 396080 17320
rect 352708 17280 352714 17292
rect 396074 17280 396080 17292
rect 396132 17280 396138 17332
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 73154 17252 73160 17264
rect 17920 17224 73160 17252
rect 17920 17212 17926 17224
rect 73154 17212 73160 17224
rect 73212 17212 73218 17264
rect 78582 17212 78588 17264
rect 78640 17252 78646 17264
rect 146938 17252 146944 17264
rect 78640 17224 146944 17252
rect 78640 17212 78646 17224
rect 146938 17212 146944 17224
rect 146996 17212 147002 17264
rect 260742 17212 260748 17264
rect 260800 17252 260806 17264
rect 489914 17252 489920 17264
rect 260800 17224 489920 17252
rect 260800 17212 260806 17224
rect 489914 17212 489920 17224
rect 489972 17212 489978 17264
rect 1104 16816 582820 16912
rect 1104 16272 582820 16368
rect 250990 15852 250996 15904
rect 251048 15892 251054 15904
rect 455690 15892 455696 15904
rect 251048 15864 455696 15892
rect 251048 15852 251054 15864
rect 455690 15852 455696 15864
rect 455748 15852 455754 15904
rect 1104 15728 582820 15824
rect 1104 15184 582820 15280
rect 1104 14640 582820 14736
rect 139302 14560 139308 14612
rect 139360 14600 139366 14612
rect 287698 14600 287704 14612
rect 139360 14572 287704 14600
rect 139360 14560 139366 14572
rect 287698 14560 287704 14572
rect 287756 14560 287762 14612
rect 84102 14492 84108 14544
rect 84160 14532 84166 14544
rect 89806 14532 89812 14544
rect 84160 14504 89812 14532
rect 84160 14492 84166 14504
rect 89806 14492 89812 14504
rect 89864 14492 89870 14544
rect 186958 14492 186964 14544
rect 187016 14532 187022 14544
rect 196802 14532 196808 14544
rect 187016 14504 196808 14532
rect 187016 14492 187022 14504
rect 196802 14492 196808 14504
rect 196860 14492 196866 14544
rect 234522 14492 234528 14544
rect 234580 14532 234586 14544
rect 390554 14532 390560 14544
rect 234580 14504 390560 14532
rect 234580 14492 234586 14504
rect 390554 14492 390560 14504
rect 390612 14492 390618 14544
rect 41322 14424 41328 14476
rect 41380 14464 41386 14476
rect 78674 14464 78680 14476
rect 41380 14436 78680 14464
rect 41380 14424 41386 14436
rect 78674 14424 78680 14436
rect 78732 14424 78738 14476
rect 85482 14424 85488 14476
rect 85540 14464 85546 14476
rect 119338 14464 119344 14476
rect 85540 14436 119344 14464
rect 85540 14424 85546 14436
rect 119338 14424 119344 14436
rect 119396 14424 119402 14476
rect 119890 14424 119896 14476
rect 119948 14464 119954 14476
rect 129734 14464 129740 14476
rect 119948 14436 129740 14464
rect 119948 14424 119954 14436
rect 129734 14424 129740 14436
rect 129792 14424 129798 14476
rect 136542 14424 136548 14476
rect 136600 14464 136606 14476
rect 168374 14464 168380 14476
rect 136600 14436 168380 14464
rect 136600 14424 136606 14436
rect 168374 14424 168380 14436
rect 168432 14424 168438 14476
rect 195238 14424 195244 14476
rect 195296 14464 195302 14476
rect 218054 14464 218060 14476
rect 195296 14436 218060 14464
rect 195296 14424 195302 14436
rect 218054 14424 218060 14436
rect 218112 14424 218118 14476
rect 258718 14424 258724 14476
rect 258776 14464 258782 14476
rect 480346 14464 480352 14476
rect 258776 14436 480352 14464
rect 258776 14424 258782 14436
rect 480346 14424 480352 14436
rect 480404 14424 480410 14476
rect 1104 14096 582820 14192
rect 1104 13552 582820 13648
rect 398098 13404 398104 13456
rect 398156 13444 398162 13456
rect 400122 13444 400128 13456
rect 398156 13416 400128 13444
rect 398156 13404 398162 13416
rect 400122 13404 400128 13416
rect 400180 13404 400186 13456
rect 240778 13132 240784 13184
rect 240836 13172 240842 13184
rect 409598 13172 409604 13184
rect 240836 13144 409604 13172
rect 240836 13132 240842 13144
rect 409598 13132 409604 13144
rect 409656 13132 409662 13184
rect 1104 13008 582820 13104
rect 1104 12464 582820 12560
rect 206922 12384 206928 12436
rect 206980 12424 206986 12436
rect 418154 12424 418160 12436
rect 206980 12396 418160 12424
rect 206980 12384 206986 12396
rect 418154 12384 418160 12396
rect 418212 12384 418218 12436
rect 202598 12316 202604 12368
rect 202656 12356 202662 12368
rect 416866 12356 416872 12368
rect 202656 12328 416872 12356
rect 202656 12316 202662 12328
rect 416866 12316 416872 12328
rect 416924 12316 416930 12368
rect 199838 12248 199844 12300
rect 199896 12288 199902 12300
rect 416774 12288 416780 12300
rect 199896 12260 416780 12288
rect 199896 12248 199902 12260
rect 416774 12248 416780 12260
rect 416832 12248 416838 12300
rect 195606 12180 195612 12232
rect 195664 12220 195670 12232
rect 415394 12220 415400 12232
rect 195664 12192 415400 12220
rect 195664 12180 195670 12192
rect 415394 12180 415400 12192
rect 415452 12180 415458 12232
rect 193030 12112 193036 12164
rect 193088 12152 193094 12164
rect 414106 12152 414112 12164
rect 193088 12124 414112 12152
rect 193088 12112 193094 12124
rect 414106 12112 414112 12124
rect 414164 12112 414170 12164
rect 188522 12044 188528 12096
rect 188580 12084 188586 12096
rect 414014 12084 414020 12096
rect 188580 12056 414020 12084
rect 188580 12044 188586 12056
rect 414014 12044 414020 12056
rect 414072 12044 414078 12096
rect 1104 11920 582820 12016
rect 186130 11840 186136 11892
rect 186188 11880 186194 11892
rect 412634 11880 412640 11892
rect 186188 11852 412640 11880
rect 186188 11840 186194 11852
rect 412634 11840 412640 11852
rect 412692 11840 412698 11892
rect 73062 11772 73068 11824
rect 73120 11812 73126 11824
rect 87046 11812 87052 11824
rect 73120 11784 87052 11812
rect 73120 11772 73126 11784
rect 87046 11772 87052 11784
rect 87104 11772 87110 11824
rect 106182 11772 106188 11824
rect 106240 11812 106246 11824
rect 125594 11812 125600 11824
rect 106240 11784 125600 11812
rect 106240 11772 106246 11784
rect 125594 11772 125600 11784
rect 125652 11772 125658 11824
rect 135438 11772 135444 11824
rect 135496 11812 135502 11824
rect 400214 11812 400220 11824
rect 135496 11784 400220 11812
rect 135496 11772 135502 11784
rect 400214 11772 400220 11784
rect 400272 11772 400278 11824
rect 60642 11704 60648 11756
rect 60700 11744 60706 11756
rect 112438 11744 112444 11756
rect 60700 11716 112444 11744
rect 60700 11704 60706 11716
rect 112438 11704 112444 11716
rect 112496 11704 112502 11756
rect 131758 11704 131764 11756
rect 131816 11744 131822 11756
rect 398926 11744 398932 11756
rect 131816 11716 398932 11744
rect 131816 11704 131822 11716
rect 398926 11704 398932 11716
rect 398984 11704 398990 11756
rect 489914 11704 489920 11756
rect 489972 11744 489978 11756
rect 491110 11744 491116 11756
rect 489972 11716 491116 11744
rect 489972 11704 489978 11716
rect 491110 11704 491116 11716
rect 491168 11704 491174 11756
rect 91002 11636 91008 11688
rect 91060 11676 91066 11688
rect 92474 11676 92480 11688
rect 91060 11648 92480 11676
rect 91060 11636 91066 11648
rect 92474 11636 92480 11648
rect 92532 11636 92538 11688
rect 211062 11636 211068 11688
rect 211120 11676 211126 11688
rect 419534 11676 419540 11688
rect 211120 11648 419540 11676
rect 211120 11636 211126 11648
rect 419534 11636 419540 11648
rect 419592 11636 419598 11688
rect 213822 11568 213828 11620
rect 213880 11608 213886 11620
rect 419626 11608 419632 11620
rect 213880 11580 419632 11608
rect 213880 11568 213886 11580
rect 419626 11568 419632 11580
rect 419684 11568 419690 11620
rect 217962 11500 217968 11552
rect 218020 11540 218026 11552
rect 420914 11540 420920 11552
rect 218020 11512 420920 11540
rect 218020 11500 218026 11512
rect 420914 11500 420920 11512
rect 420972 11500 420978 11552
rect 1104 11376 582820 11472
rect 220446 11296 220452 11348
rect 220504 11336 220510 11348
rect 422386 11336 422392 11348
rect 220504 11308 422392 11336
rect 220504 11296 220510 11308
rect 422386 11296 422392 11308
rect 422444 11296 422450 11348
rect 224770 11228 224776 11280
rect 224828 11268 224834 11280
rect 422294 11268 422300 11280
rect 224828 11240 422300 11268
rect 224828 11228 224834 11240
rect 422294 11228 422300 11240
rect 422352 11228 422358 11280
rect 227438 11160 227444 11212
rect 227496 11200 227502 11212
rect 423674 11200 423680 11212
rect 227496 11172 423680 11200
rect 227496 11160 227502 11172
rect 423674 11160 423680 11172
rect 423732 11160 423738 11212
rect 238662 11092 238668 11144
rect 238720 11132 238726 11144
rect 292298 11132 292304 11144
rect 238720 11104 292304 11132
rect 238720 11092 238726 11104
rect 292298 11092 292304 11104
rect 292356 11092 292362 11144
rect 292408 11104 292712 11132
rect 270034 11024 270040 11076
rect 270092 11064 270098 11076
rect 282638 11064 282644 11076
rect 270092 11036 282644 11064
rect 270092 11024 270098 11036
rect 282638 11024 282644 11036
rect 282696 11024 282702 11076
rect 292408 11064 292436 11104
rect 282748 11036 292436 11064
rect 292485 11067 292543 11073
rect 181990 10956 181996 11008
rect 182048 10996 182054 11008
rect 282748 10996 282776 11036
rect 292485 11033 292497 11067
rect 292531 11064 292543 11067
rect 292574 11064 292580 11076
rect 292531 11036 292580 11064
rect 292531 11033 292543 11036
rect 292485 11027 292543 11033
rect 292574 11024 292580 11036
rect 292632 11024 292638 11076
rect 292684 11064 292712 11104
rect 292942 11092 292948 11144
rect 293000 11132 293006 11144
rect 426434 11132 426440 11144
rect 293000 11104 426440 11132
rect 293000 11092 293006 11104
rect 426434 11092 426440 11104
rect 426492 11092 426498 11144
rect 292684 11036 302372 11064
rect 182048 10968 282776 10996
rect 282825 10999 282883 11005
rect 182048 10956 182054 10968
rect 282825 10965 282837 10999
rect 282871 10996 282883 10999
rect 292301 10999 292359 11005
rect 292301 10996 292313 10999
rect 282871 10968 292313 10996
rect 282871 10965 282883 10968
rect 282825 10959 282883 10965
rect 292301 10965 292313 10968
rect 292347 10965 292359 10999
rect 292301 10959 292359 10965
rect 292393 10999 292451 11005
rect 292393 10965 292405 10999
rect 292439 10996 292451 10999
rect 302237 10999 302295 11005
rect 302237 10996 302249 10999
rect 292439 10968 302249 10996
rect 292439 10965 292451 10968
rect 292393 10959 292451 10965
rect 302237 10965 302249 10968
rect 302283 10965 302295 10999
rect 302344 10996 302372 11036
rect 302510 11024 302516 11076
rect 302568 11064 302574 11076
rect 434714 11064 434720 11076
rect 302568 11036 434720 11064
rect 302568 11024 302574 11036
rect 434714 11024 434720 11036
rect 434772 11024 434778 11076
rect 411346 10996 411352 11008
rect 302344 10968 411352 10996
rect 302237 10959 302295 10965
rect 411346 10956 411352 10968
rect 411404 10956 411410 11008
rect 1104 10832 582820 10928
rect 177850 10752 177856 10804
rect 177908 10792 177914 10804
rect 277581 10795 277639 10801
rect 277581 10792 277593 10795
rect 177908 10764 277593 10792
rect 177908 10752 177914 10764
rect 277581 10761 277593 10764
rect 277627 10761 277639 10795
rect 286873 10795 286931 10801
rect 286873 10792 286885 10795
rect 277581 10755 277639 10761
rect 277688 10764 286885 10792
rect 175182 10684 175188 10736
rect 175240 10724 175246 10736
rect 277688 10724 277716 10764
rect 286873 10761 286885 10764
rect 286919 10761 286931 10795
rect 302237 10795 302295 10801
rect 302237 10792 302249 10795
rect 286873 10755 286931 10761
rect 286980 10764 302249 10792
rect 286980 10724 287008 10764
rect 302237 10761 302249 10764
rect 302283 10761 302295 10795
rect 302237 10755 302295 10761
rect 302326 10752 302332 10804
rect 302384 10792 302390 10804
rect 411254 10792 411260 10804
rect 302384 10764 411260 10792
rect 302384 10752 302390 10764
rect 411254 10752 411260 10764
rect 411312 10752 411318 10804
rect 307205 10727 307263 10733
rect 175240 10696 277716 10724
rect 277780 10696 287008 10724
rect 287072 10696 307156 10724
rect 175240 10684 175246 10696
rect 170766 10616 170772 10668
rect 170824 10656 170830 10668
rect 277780 10656 277808 10696
rect 287072 10656 287100 10696
rect 307128 10656 307156 10696
rect 307205 10693 307217 10727
rect 307251 10724 307263 10727
rect 307251 10696 311756 10724
rect 307251 10693 307263 10696
rect 307205 10687 307263 10693
rect 311621 10659 311679 10665
rect 311621 10656 311633 10659
rect 170824 10628 277808 10656
rect 277872 10628 287100 10656
rect 287164 10628 307064 10656
rect 307128 10628 311633 10656
rect 170824 10616 170830 10628
rect 168282 10548 168288 10600
rect 168340 10588 168346 10600
rect 277872 10588 277900 10628
rect 287164 10588 287192 10628
rect 168340 10560 277900 10588
rect 277964 10560 287192 10588
rect 287241 10591 287299 10597
rect 168340 10548 168346 10560
rect 163682 10480 163688 10532
rect 163740 10520 163746 10532
rect 277964 10520 277992 10560
rect 287241 10557 287253 10591
rect 287287 10588 287299 10591
rect 287609 10591 287667 10597
rect 287609 10588 287621 10591
rect 287287 10560 287621 10588
rect 287287 10557 287299 10560
rect 287241 10551 287299 10557
rect 287609 10557 287621 10560
rect 287655 10557 287667 10591
rect 306377 10591 306435 10597
rect 287609 10551 287667 10557
rect 287716 10560 306328 10588
rect 287716 10520 287744 10560
rect 163740 10492 277992 10520
rect 278056 10492 287744 10520
rect 287793 10523 287851 10529
rect 163740 10480 163746 10492
rect 128170 10412 128176 10464
rect 128228 10452 128234 10464
rect 278056 10452 278084 10492
rect 287793 10489 287805 10523
rect 287839 10520 287851 10523
rect 292301 10523 292359 10529
rect 292301 10520 292313 10523
rect 287839 10492 292313 10520
rect 287839 10489 287851 10492
rect 287793 10483 287851 10489
rect 292301 10489 292313 10492
rect 292347 10489 292359 10523
rect 292301 10483 292359 10489
rect 292390 10480 292396 10532
rect 292448 10520 292454 10532
rect 302326 10520 302332 10532
rect 292448 10492 302332 10520
rect 292448 10480 292454 10492
rect 302326 10480 302332 10492
rect 302384 10480 302390 10532
rect 302421 10523 302479 10529
rect 302421 10489 302433 10523
rect 302467 10520 302479 10523
rect 306193 10523 306251 10529
rect 306193 10520 306205 10523
rect 302467 10492 306205 10520
rect 302467 10489 302479 10492
rect 302421 10483 302479 10489
rect 306193 10489 306205 10492
rect 306239 10489 306251 10523
rect 306300 10520 306328 10560
rect 306377 10557 306389 10591
rect 306423 10588 306435 10591
rect 306929 10591 306987 10597
rect 306929 10588 306941 10591
rect 306423 10560 306941 10588
rect 306423 10557 306435 10560
rect 306377 10551 306435 10557
rect 306929 10557 306941 10560
rect 306975 10557 306987 10591
rect 307036 10588 307064 10628
rect 311621 10625 311633 10628
rect 311667 10625 311679 10659
rect 311728 10656 311756 10696
rect 311802 10684 311808 10736
rect 311860 10724 311866 10736
rect 409874 10724 409880 10736
rect 311860 10696 409880 10724
rect 311860 10684 311866 10696
rect 409874 10684 409880 10696
rect 409932 10684 409938 10736
rect 408494 10656 408500 10668
rect 311728 10628 408500 10656
rect 311621 10619 311679 10625
rect 408494 10616 408500 10628
rect 408552 10616 408558 10668
rect 311529 10591 311587 10597
rect 311529 10588 311541 10591
rect 307036 10560 311541 10588
rect 306929 10551 306987 10557
rect 311529 10557 311541 10560
rect 311575 10557 311587 10591
rect 311529 10551 311587 10557
rect 311897 10591 311955 10597
rect 311897 10557 311909 10591
rect 311943 10588 311955 10591
rect 408586 10588 408592 10600
rect 311943 10560 408592 10588
rect 311943 10557 311955 10560
rect 311897 10551 311955 10557
rect 408586 10548 408592 10560
rect 408644 10548 408650 10600
rect 311805 10523 311863 10529
rect 306300 10492 311756 10520
rect 306193 10483 306251 10489
rect 128228 10424 278084 10452
rect 278133 10455 278191 10461
rect 128228 10412 128234 10424
rect 278133 10421 278145 10455
rect 278179 10452 278191 10455
rect 282733 10455 282791 10461
rect 282733 10452 282745 10455
rect 278179 10424 282745 10452
rect 278179 10421 278191 10424
rect 278133 10415 278191 10421
rect 282733 10421 282745 10424
rect 282779 10421 282791 10455
rect 282733 10415 282791 10421
rect 282822 10412 282828 10464
rect 282880 10452 282886 10464
rect 311526 10452 311532 10464
rect 282880 10424 311532 10452
rect 282880 10412 282886 10424
rect 311526 10412 311532 10424
rect 311584 10412 311590 10464
rect 311728 10452 311756 10492
rect 311805 10489 311817 10523
rect 311851 10520 311863 10523
rect 407114 10520 407120 10532
rect 311851 10492 407120 10520
rect 311851 10489 311863 10492
rect 311805 10483 311863 10489
rect 407114 10480 407120 10492
rect 407172 10480 407178 10532
rect 398834 10452 398840 10464
rect 311728 10424 398840 10452
rect 398834 10412 398840 10424
rect 398892 10412 398898 10464
rect 1104 10288 582820 10384
rect 252370 10208 252376 10260
rect 252428 10248 252434 10260
rect 311434 10248 311440 10260
rect 252428 10220 311440 10248
rect 252428 10208 252434 10220
rect 311434 10208 311440 10220
rect 311492 10208 311498 10260
rect 311802 10208 311808 10260
rect 311860 10248 311866 10260
rect 320174 10248 320180 10260
rect 311860 10220 320180 10248
rect 311860 10208 311866 10220
rect 320174 10208 320180 10220
rect 320232 10208 320238 10260
rect 372522 10208 372528 10260
rect 372580 10248 372586 10260
rect 477586 10248 477592 10260
rect 372580 10220 477592 10248
rect 372580 10208 372586 10220
rect 477586 10208 477592 10220
rect 477644 10208 477650 10260
rect 255222 10140 255228 10192
rect 255280 10180 255286 10192
rect 302237 10183 302295 10189
rect 302237 10180 302249 10183
rect 255280 10152 302249 10180
rect 255280 10140 255286 10152
rect 302237 10149 302249 10152
rect 302283 10149 302295 10183
rect 302237 10143 302295 10149
rect 302329 10183 302387 10189
rect 302329 10149 302341 10183
rect 302375 10180 302387 10183
rect 307205 10183 307263 10189
rect 307205 10180 307217 10183
rect 302375 10152 307217 10180
rect 302375 10149 302387 10152
rect 302329 10143 302387 10149
rect 307205 10149 307217 10152
rect 307251 10149 307263 10183
rect 307205 10143 307263 10149
rect 307297 10183 307355 10189
rect 307297 10149 307309 10183
rect 307343 10180 307355 10183
rect 311618 10180 311624 10192
rect 307343 10152 311624 10180
rect 307343 10149 307355 10152
rect 307297 10143 307355 10149
rect 311618 10140 311624 10152
rect 311676 10140 311682 10192
rect 311710 10140 311716 10192
rect 311768 10180 311774 10192
rect 321646 10180 321652 10192
rect 311768 10152 321652 10180
rect 311768 10140 311774 10152
rect 321646 10140 321652 10152
rect 321704 10140 321710 10192
rect 372430 10140 372436 10192
rect 372488 10180 372494 10192
rect 474550 10180 474556 10192
rect 372488 10152 474556 10180
rect 372488 10140 372494 10152
rect 474550 10140 474556 10152
rect 474608 10140 474614 10192
rect 259362 10072 259368 10124
rect 259420 10112 259426 10124
rect 316126 10112 316132 10124
rect 259420 10084 316132 10112
rect 259420 10072 259426 10084
rect 316126 10072 316132 10084
rect 316184 10072 316190 10124
rect 369670 10072 369676 10124
rect 369728 10112 369734 10124
rect 467466 10112 467472 10124
rect 369728 10084 467472 10112
rect 369728 10072 369734 10084
rect 467466 10072 467472 10084
rect 467524 10072 467530 10124
rect 261754 10004 261760 10056
rect 261812 10044 261818 10056
rect 307113 10047 307171 10053
rect 261812 10016 307064 10044
rect 261812 10004 261818 10016
rect 266078 9936 266084 9988
rect 266136 9976 266142 9988
rect 306929 9979 306987 9985
rect 306929 9976 306941 9979
rect 266136 9948 306941 9976
rect 266136 9936 266142 9948
rect 306929 9945 306941 9948
rect 306975 9945 306987 9979
rect 307036 9976 307064 10016
rect 307113 10013 307125 10047
rect 307159 10044 307171 10047
rect 317414 10044 317420 10056
rect 307159 10016 317420 10044
rect 307159 10013 307171 10016
rect 307113 10007 307171 10013
rect 317414 10004 317420 10016
rect 317472 10004 317478 10056
rect 316034 9976 316040 9988
rect 307036 9948 316040 9976
rect 306929 9939 306987 9945
rect 316034 9936 316040 9948
rect 316092 9936 316098 9988
rect 268838 9868 268844 9920
rect 268896 9908 268902 9920
rect 318794 9908 318800 9920
rect 268896 9880 318800 9908
rect 268896 9868 268902 9880
rect 318794 9868 318800 9880
rect 318852 9868 318858 9920
rect 1104 9744 582820 9840
rect 273070 9664 273076 9716
rect 273128 9704 273134 9716
rect 318886 9704 318892 9716
rect 273128 9676 318892 9704
rect 273128 9664 273134 9676
rect 318886 9664 318892 9676
rect 318944 9664 318950 9716
rect 190822 9596 190828 9648
rect 190880 9636 190886 9648
rect 298094 9636 298100 9648
rect 190880 9608 298100 9636
rect 190880 9596 190886 9608
rect 298094 9596 298100 9608
rect 298152 9596 298158 9648
rect 302237 9639 302295 9645
rect 302237 9605 302249 9639
rect 302283 9636 302295 9639
rect 314654 9636 314660 9648
rect 302283 9608 314660 9636
rect 302283 9605 302295 9608
rect 302237 9599 302295 9605
rect 314654 9596 314660 9608
rect 314712 9596 314718 9648
rect 361482 9596 361488 9648
rect 361540 9636 361546 9648
rect 432046 9636 432052 9648
rect 361540 9608 432052 9636
rect 361540 9596 361546 9608
rect 432046 9596 432052 9608
rect 432104 9596 432110 9648
rect 187326 9528 187332 9580
rect 187384 9568 187390 9580
rect 296714 9568 296720 9580
rect 187384 9540 296720 9568
rect 187384 9528 187390 9540
rect 296714 9528 296720 9540
rect 296772 9528 296778 9580
rect 362862 9528 362868 9580
rect 362920 9568 362926 9580
rect 435542 9568 435548 9580
rect 362920 9540 435548 9568
rect 362920 9528 362926 9540
rect 435542 9528 435548 9540
rect 435600 9528 435606 9580
rect 183738 9460 183744 9512
rect 183796 9500 183802 9512
rect 284113 9503 284171 9509
rect 284113 9500 284125 9503
rect 183796 9472 284125 9500
rect 183796 9460 183802 9472
rect 284113 9469 284125 9472
rect 284159 9469 284171 9503
rect 292390 9500 292396 9512
rect 284113 9463 284171 9469
rect 284220 9472 292396 9500
rect 180242 9392 180248 9444
rect 180300 9432 180306 9444
rect 284220 9432 284248 9472
rect 292390 9460 292396 9472
rect 292448 9460 292454 9512
rect 292485 9503 292543 9509
rect 292485 9469 292497 9503
rect 292531 9500 292543 9503
rect 293954 9500 293960 9512
rect 292531 9472 293960 9500
rect 292531 9469 292543 9472
rect 292485 9463 292543 9469
rect 293954 9460 293960 9472
rect 294012 9460 294018 9512
rect 362770 9460 362776 9512
rect 362828 9500 362834 9512
rect 439130 9500 439136 9512
rect 362828 9472 439136 9500
rect 362828 9460 362834 9472
rect 439130 9460 439136 9472
rect 439188 9460 439194 9512
rect 294046 9432 294052 9444
rect 180300 9404 284248 9432
rect 284312 9404 294052 9432
rect 180300 9392 180306 9404
rect 176654 9324 176660 9376
rect 176712 9364 176718 9376
rect 284312 9364 284340 9404
rect 294046 9392 294052 9404
rect 294104 9392 294110 9444
rect 364242 9392 364248 9444
rect 364300 9432 364306 9444
rect 442626 9432 442632 9444
rect 364300 9404 442632 9432
rect 364300 9392 364306 9404
rect 442626 9392 442632 9404
rect 442684 9392 442690 9444
rect 176712 9336 284340 9364
rect 284389 9367 284447 9373
rect 176712 9324 176718 9336
rect 284389 9333 284401 9367
rect 284435 9364 284447 9367
rect 287517 9367 287575 9373
rect 287517 9364 287529 9367
rect 284435 9336 287529 9364
rect 284435 9333 284447 9336
rect 284389 9327 284447 9333
rect 287517 9333 287529 9336
rect 287563 9333 287575 9367
rect 287517 9327 287575 9333
rect 287609 9367 287667 9373
rect 287609 9333 287621 9367
rect 287655 9364 287667 9367
rect 292666 9364 292672 9376
rect 287655 9336 292672 9364
rect 287655 9333 287667 9336
rect 287609 9327 287667 9333
rect 292666 9324 292672 9336
rect 292724 9324 292730 9376
rect 292942 9324 292948 9376
rect 293000 9364 293006 9376
rect 295334 9364 295340 9376
rect 293000 9336 295340 9364
rect 293000 9324 293006 9336
rect 295334 9324 295340 9336
rect 295392 9324 295398 9376
rect 365530 9324 365536 9376
rect 365588 9364 365594 9376
rect 446214 9364 446220 9376
rect 365588 9336 446220 9364
rect 365588 9324 365594 9336
rect 446214 9324 446220 9336
rect 446272 9324 446278 9376
rect 1104 9200 582820 9296
rect 173158 9120 173164 9172
rect 173216 9160 173222 9172
rect 292301 9163 292359 9169
rect 292301 9160 292313 9163
rect 173216 9132 292313 9160
rect 173216 9120 173222 9132
rect 292301 9129 292313 9132
rect 292347 9129 292359 9163
rect 292301 9123 292359 9129
rect 292485 9163 292543 9169
rect 292485 9129 292497 9163
rect 292531 9160 292543 9163
rect 296990 9160 296996 9172
rect 292531 9132 296996 9160
rect 292531 9129 292543 9132
rect 292485 9123 292543 9129
rect 296990 9120 296996 9132
rect 297048 9120 297054 9172
rect 366910 9120 366916 9172
rect 366968 9160 366974 9172
rect 366968 9132 373856 9160
rect 366968 9120 366974 9132
rect 169570 9052 169576 9104
rect 169628 9092 169634 9104
rect 287609 9095 287667 9101
rect 287609 9092 287621 9095
rect 169628 9064 287621 9092
rect 169628 9052 169634 9064
rect 287609 9061 287621 9064
rect 287655 9061 287667 9095
rect 292850 9092 292856 9104
rect 287609 9055 287667 9061
rect 287716 9064 292856 9092
rect 66714 8984 66720 9036
rect 66772 9024 66778 9036
rect 115198 9024 115204 9036
rect 66772 8996 115204 9024
rect 66772 8984 66778 8996
rect 115198 8984 115204 8996
rect 115256 8984 115262 9036
rect 166074 8984 166080 9036
rect 166132 9024 166138 9036
rect 287716 9024 287744 9064
rect 292850 9052 292856 9064
rect 292908 9052 292914 9104
rect 365622 9052 365628 9104
rect 365680 9092 365686 9104
rect 369670 9092 369676 9104
rect 365680 9064 369676 9092
rect 365680 9052 365686 9064
rect 369670 9052 369676 9064
rect 369728 9052 369734 9104
rect 369762 9052 369768 9104
rect 369820 9092 369826 9104
rect 373718 9092 373724 9104
rect 369820 9064 373724 9092
rect 369820 9052 369826 9064
rect 373718 9052 373724 9064
rect 373776 9052 373782 9104
rect 373828 9092 373856 9132
rect 373902 9120 373908 9172
rect 373960 9160 373966 9172
rect 449802 9160 449808 9172
rect 373960 9132 449808 9160
rect 373960 9120 373966 9132
rect 449802 9120 449808 9132
rect 449860 9120 449866 9172
rect 456886 9092 456892 9104
rect 373828 9064 456892 9092
rect 456886 9052 456892 9064
rect 456944 9052 456950 9104
rect 166132 8996 287744 9024
rect 287793 9027 287851 9033
rect 166132 8984 166138 8996
rect 287793 8993 287805 9027
rect 287839 9024 287851 9027
rect 292393 9027 292451 9033
rect 292393 9024 292405 9027
rect 287839 8996 292405 9024
rect 287839 8993 287851 8996
rect 287793 8987 287851 8993
rect 292393 8993 292405 8996
rect 292439 8993 292451 9027
rect 292393 8987 292451 8993
rect 292485 9027 292543 9033
rect 292485 8993 292497 9027
rect 292531 9024 292543 9027
rect 321554 9024 321560 9036
rect 292531 8996 321560 9024
rect 292531 8993 292543 8996
rect 292485 8987 292543 8993
rect 321554 8984 321560 8996
rect 321612 8984 321618 9036
rect 368382 8984 368388 9036
rect 368440 9024 368446 9036
rect 460382 9024 460388 9036
rect 368440 8996 460388 9024
rect 368440 8984 368446 8996
rect 460382 8984 460388 8996
rect 460440 8984 460446 9036
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 74534 8956 74540 8968
rect 21876 8928 74540 8956
rect 21876 8916 21882 8928
rect 74534 8916 74540 8928
rect 74592 8916 74598 8968
rect 79686 8916 79692 8968
rect 79744 8956 79750 8968
rect 89714 8956 89720 8968
rect 79744 8928 89720 8956
rect 79744 8916 79750 8928
rect 89714 8916 89720 8928
rect 89772 8916 89778 8968
rect 102226 8916 102232 8968
rect 102284 8956 102290 8968
rect 124306 8956 124312 8968
rect 102284 8928 124312 8956
rect 102284 8916 102290 8928
rect 124306 8916 124312 8928
rect 124364 8916 124370 8968
rect 130562 8916 130568 8968
rect 130620 8956 130626 8968
rect 273254 8956 273260 8968
rect 130620 8928 273260 8956
rect 130620 8916 130626 8928
rect 273254 8916 273260 8928
rect 273312 8916 273318 8968
rect 273346 8916 273352 8968
rect 273404 8956 273410 8968
rect 305086 8956 305092 8968
rect 273404 8928 305092 8956
rect 273404 8916 273410 8928
rect 305086 8916 305092 8928
rect 305144 8916 305150 8968
rect 354490 8916 354496 8968
rect 354548 8956 354554 8968
rect 393314 8956 393320 8968
rect 354548 8928 393320 8956
rect 354548 8916 354554 8928
rect 393314 8916 393320 8928
rect 393372 8916 393378 8968
rect 393406 8916 393412 8968
rect 393464 8956 393470 8968
rect 463970 8956 463976 8968
rect 393464 8928 463976 8956
rect 393464 8916 393470 8928
rect 463970 8916 463976 8928
rect 464028 8916 464034 8968
rect 194410 8848 194416 8900
rect 194468 8888 194474 8900
rect 299566 8888 299572 8900
rect 194468 8860 299572 8888
rect 194468 8848 194474 8860
rect 299566 8848 299572 8860
rect 299624 8848 299630 8900
rect 360102 8848 360108 8900
rect 360160 8888 360166 8900
rect 428458 8888 428464 8900
rect 360160 8860 428464 8888
rect 360160 8848 360166 8860
rect 428458 8848 428464 8860
rect 428516 8848 428522 8900
rect 197906 8780 197912 8832
rect 197964 8820 197970 8832
rect 299474 8820 299480 8832
rect 197964 8792 299480 8820
rect 197964 8780 197970 8792
rect 299474 8780 299480 8792
rect 299532 8780 299538 8832
rect 360010 8780 360016 8832
rect 360068 8820 360074 8832
rect 424962 8820 424968 8832
rect 360068 8792 424968 8820
rect 360068 8780 360074 8792
rect 424962 8780 424968 8792
rect 425020 8780 425026 8832
rect 1104 8656 582820 8752
rect 201494 8576 201500 8628
rect 201552 8616 201558 8628
rect 300854 8616 300860 8628
rect 201552 8588 300860 8616
rect 201552 8576 201558 8588
rect 300854 8576 300860 8588
rect 300912 8576 300918 8628
rect 358722 8576 358728 8628
rect 358780 8616 358786 8628
rect 421374 8616 421380 8628
rect 358780 8588 421380 8616
rect 358780 8576 358786 8588
rect 421374 8576 421380 8588
rect 421432 8576 421438 8628
rect 205082 8508 205088 8560
rect 205140 8548 205146 8560
rect 302234 8548 302240 8560
rect 205140 8520 302240 8548
rect 205140 8508 205146 8520
rect 302234 8508 302240 8520
rect 302292 8508 302298 8560
rect 357342 8508 357348 8560
rect 357400 8548 357406 8560
rect 417878 8548 417884 8560
rect 357400 8520 417884 8548
rect 357400 8508 357406 8520
rect 417878 8508 417884 8520
rect 417936 8508 417942 8560
rect 208578 8440 208584 8492
rect 208636 8480 208642 8492
rect 302418 8480 302424 8492
rect 208636 8452 302424 8480
rect 208636 8440 208642 8452
rect 302418 8440 302424 8452
rect 302476 8440 302482 8492
rect 357250 8440 357256 8492
rect 357308 8480 357314 8492
rect 414290 8480 414296 8492
rect 357308 8452 414296 8480
rect 357308 8440 357314 8452
rect 414290 8440 414296 8452
rect 414348 8440 414354 8492
rect 212166 8372 212172 8424
rect 212224 8412 212230 8424
rect 303614 8412 303620 8424
rect 212224 8384 303620 8412
rect 212224 8372 212230 8384
rect 303614 8372 303620 8384
rect 303672 8372 303678 8424
rect 355962 8372 355968 8424
rect 356020 8412 356026 8424
rect 410794 8412 410800 8424
rect 356020 8384 410800 8412
rect 356020 8372 356026 8384
rect 410794 8372 410800 8384
rect 410852 8372 410858 8424
rect 215662 8304 215668 8356
rect 215720 8344 215726 8356
rect 304994 8344 305000 8356
rect 215720 8316 305000 8344
rect 215720 8304 215726 8316
rect 304994 8304 305000 8316
rect 305052 8304 305058 8356
rect 354582 8304 354588 8356
rect 354640 8344 354646 8356
rect 407206 8344 407212 8356
rect 354640 8316 407212 8344
rect 354640 8304 354646 8316
rect 407206 8304 407212 8316
rect 407264 8304 407270 8356
rect 219250 8236 219256 8288
rect 219308 8276 219314 8288
rect 248874 8276 248880 8288
rect 219308 8248 248880 8276
rect 219308 8236 219314 8248
rect 248874 8236 248880 8248
rect 248932 8236 248938 8288
rect 253201 8279 253259 8285
rect 253201 8245 253213 8279
rect 253247 8276 253259 8279
rect 430850 8276 430856 8288
rect 253247 8248 430856 8276
rect 253247 8245 253259 8248
rect 253201 8239 253259 8245
rect 430850 8236 430856 8248
rect 430908 8236 430914 8288
rect 1104 8112 582820 8208
rect 245562 8032 245568 8084
rect 245620 8072 245626 8084
rect 253201 8075 253259 8081
rect 253201 8072 253213 8075
rect 245620 8044 253213 8072
rect 245620 8032 245626 8044
rect 253201 8041 253213 8044
rect 253247 8041 253259 8075
rect 253201 8035 253259 8041
rect 253293 8075 253351 8081
rect 253293 8041 253305 8075
rect 253339 8072 253351 8075
rect 434438 8072 434444 8084
rect 253339 8044 434444 8072
rect 253339 8041 253351 8044
rect 253293 8035 253351 8041
rect 434438 8032 434444 8044
rect 434496 8032 434502 8084
rect 246942 7964 246948 8016
rect 247000 8004 247006 8016
rect 437934 8004 437940 8016
rect 247000 7976 437940 8004
rect 247000 7964 247006 7976
rect 437934 7964 437940 7976
rect 437992 7964 437998 8016
rect 248322 7896 248328 7948
rect 248380 7936 248386 7948
rect 441522 7936 441528 7948
rect 248380 7908 441528 7936
rect 248380 7896 248386 7908
rect 441522 7896 441528 7908
rect 441580 7896 441586 7948
rect 248230 7828 248236 7880
rect 248288 7868 248294 7880
rect 445018 7868 445024 7880
rect 248288 7840 445024 7868
rect 248288 7828 248294 7840
rect 445018 7828 445024 7840
rect 445076 7828 445082 7880
rect 251082 7760 251088 7812
rect 251140 7800 251146 7812
rect 253477 7803 253535 7809
rect 251140 7772 253428 7800
rect 251140 7760 251146 7772
rect 245470 7692 245476 7744
rect 245528 7732 245534 7744
rect 253293 7735 253351 7741
rect 253293 7732 253305 7735
rect 245528 7704 253305 7732
rect 245528 7692 245534 7704
rect 253293 7701 253305 7704
rect 253339 7701 253351 7735
rect 253400 7732 253428 7772
rect 253477 7769 253489 7803
rect 253523 7800 253535 7803
rect 448606 7800 448612 7812
rect 253523 7772 448612 7800
rect 253523 7769 253535 7772
rect 253477 7763 253535 7769
rect 448606 7760 448612 7772
rect 448664 7760 448670 7812
rect 452102 7732 452108 7744
rect 253400 7704 452108 7732
rect 253293 7695 253351 7701
rect 452102 7692 452108 7704
rect 452160 7692 452166 7744
rect 1104 7568 582820 7664
rect 244182 7488 244188 7540
rect 244240 7528 244246 7540
rect 427262 7528 427268 7540
rect 244240 7500 427268 7528
rect 244240 7488 244246 7500
rect 427262 7488 427268 7500
rect 427320 7488 427326 7540
rect 463881 7531 463939 7537
rect 463881 7497 463893 7531
rect 463927 7528 463939 7531
rect 465813 7531 465871 7537
rect 465813 7528 465825 7531
rect 463927 7500 465825 7528
rect 463927 7497 463939 7500
rect 463881 7491 463939 7497
rect 465813 7497 465825 7500
rect 465859 7497 465871 7531
rect 465813 7491 465871 7497
rect 242802 7420 242808 7472
rect 242860 7460 242866 7472
rect 412634 7460 412640 7472
rect 242860 7432 412640 7460
rect 242860 7420 242866 7432
rect 412634 7420 412640 7432
rect 412692 7420 412698 7472
rect 412726 7420 412732 7472
rect 412784 7460 412790 7472
rect 577406 7460 577412 7472
rect 412784 7432 577412 7460
rect 412784 7420 412790 7432
rect 577406 7420 577412 7432
rect 577464 7420 577470 7472
rect 249702 7352 249708 7404
rect 249760 7392 249766 7404
rect 253477 7395 253535 7401
rect 253477 7392 253489 7395
rect 249760 7364 253489 7392
rect 249760 7352 249766 7364
rect 253477 7361 253489 7364
rect 253523 7361 253535 7395
rect 253477 7355 253535 7361
rect 284202 7352 284208 7404
rect 284260 7392 284266 7404
rect 292485 7395 292543 7401
rect 292485 7392 292497 7395
rect 284260 7364 292497 7392
rect 284260 7352 284266 7364
rect 292485 7361 292497 7364
rect 292531 7361 292543 7395
rect 292485 7355 292543 7361
rect 367002 7352 367008 7404
rect 367060 7392 367066 7404
rect 453298 7392 453304 7404
rect 367060 7364 453304 7392
rect 367060 7352 367066 7364
rect 453298 7352 453304 7364
rect 453356 7352 453362 7404
rect 465721 7395 465779 7401
rect 465721 7361 465733 7395
rect 465767 7392 465779 7395
rect 471054 7392 471060 7404
rect 465767 7364 471060 7392
rect 465767 7361 465779 7364
rect 465721 7355 465779 7361
rect 471054 7352 471060 7364
rect 471112 7352 471118 7404
rect 394510 7284 394516 7336
rect 394568 7324 394574 7336
rect 398650 7324 398656 7336
rect 394568 7296 398656 7324
rect 394568 7284 394574 7296
rect 398650 7284 398656 7296
rect 398708 7284 398714 7336
rect 398742 7284 398748 7336
rect 398800 7324 398806 7336
rect 400033 7327 400091 7333
rect 400033 7324 400045 7327
rect 398800 7296 400045 7324
rect 398800 7284 398806 7296
rect 400033 7293 400045 7296
rect 400079 7293 400091 7327
rect 573910 7324 573916 7336
rect 400033 7287 400091 7293
rect 400140 7296 573916 7324
rect 397362 7216 397368 7268
rect 397420 7256 397426 7268
rect 400140 7256 400168 7296
rect 573910 7284 573916 7296
rect 573968 7284 573974 7336
rect 570322 7256 570328 7268
rect 397420 7228 400168 7256
rect 400232 7228 570328 7256
rect 397420 7216 397426 7228
rect 397270 7148 397276 7200
rect 397328 7188 397334 7200
rect 400232 7188 400260 7228
rect 570322 7216 570328 7228
rect 570380 7216 570386 7268
rect 397328 7160 400260 7188
rect 400309 7191 400367 7197
rect 397328 7148 397334 7160
rect 400309 7157 400321 7191
rect 400355 7188 400367 7191
rect 408310 7188 408316 7200
rect 400355 7160 408316 7188
rect 400355 7157 400367 7160
rect 400309 7151 400367 7157
rect 408310 7148 408316 7160
rect 408368 7148 408374 7200
rect 408402 7148 408408 7200
rect 408460 7188 408466 7200
rect 566826 7188 566832 7200
rect 408460 7160 566832 7188
rect 408460 7148 408466 7160
rect 566826 7148 566832 7160
rect 566884 7148 566890 7200
rect 1104 7024 582820 7120
rect 395982 6944 395988 6996
rect 396040 6984 396046 6996
rect 398834 6984 398840 6996
rect 396040 6956 398840 6984
rect 396040 6944 396046 6956
rect 398834 6944 398840 6956
rect 398892 6944 398898 6996
rect 398926 6944 398932 6996
rect 398984 6984 398990 6996
rect 563238 6984 563244 6996
rect 398984 6956 563244 6984
rect 398984 6944 398990 6956
rect 563238 6944 563244 6956
rect 563296 6944 563302 6996
rect 371142 6876 371148 6928
rect 371200 6916 371206 6928
rect 465721 6919 465779 6925
rect 465721 6916 465733 6919
rect 371200 6888 465733 6916
rect 371200 6876 371206 6888
rect 465721 6885 465733 6888
rect 465767 6885 465779 6919
rect 465721 6879 465779 6885
rect 465813 6919 465871 6925
rect 465813 6885 465825 6919
rect 465859 6916 465871 6919
rect 502245 6919 502303 6925
rect 502245 6916 502257 6919
rect 465859 6888 502257 6916
rect 465859 6885 465871 6888
rect 465813 6879 465871 6885
rect 502245 6885 502257 6888
rect 502291 6885 502303 6919
rect 502245 6879 502303 6885
rect 293678 6808 293684 6860
rect 293736 6848 293742 6860
rect 324406 6848 324412 6860
rect 293736 6820 324412 6848
rect 293736 6808 293742 6820
rect 324406 6808 324412 6820
rect 324464 6808 324470 6860
rect 345750 6848 345756 6860
rect 335326 6820 345756 6848
rect 290182 6740 290188 6792
rect 290240 6780 290246 6792
rect 324314 6780 324320 6792
rect 290240 6752 324320 6780
rect 290240 6740 290246 6752
rect 324314 6740 324320 6752
rect 324372 6740 324378 6792
rect 325602 6740 325608 6792
rect 325660 6780 325666 6792
rect 332594 6780 332600 6792
rect 325660 6752 332600 6780
rect 325660 6740 325666 6752
rect 332594 6740 332600 6752
rect 332652 6740 332658 6792
rect 286594 6672 286600 6724
rect 286652 6712 286658 6724
rect 322934 6712 322940 6724
rect 286652 6684 322940 6712
rect 286652 6672 286658 6684
rect 322934 6672 322940 6684
rect 322992 6672 322998 6724
rect 323026 6672 323032 6724
rect 323084 6712 323090 6724
rect 331306 6712 331312 6724
rect 323084 6684 331312 6712
rect 323084 6672 323090 6684
rect 331306 6672 331312 6684
rect 331364 6672 331370 6724
rect 223482 6604 223488 6656
rect 223540 6644 223546 6656
rect 335326 6644 335354 6820
rect 345750 6808 345756 6820
rect 345808 6808 345814 6860
rect 346210 6808 346216 6860
rect 346268 6848 346274 6860
rect 375282 6848 375288 6860
rect 346268 6820 375288 6848
rect 346268 6808 346274 6820
rect 375282 6808 375288 6820
rect 375340 6808 375346 6860
rect 386230 6808 386236 6860
rect 386288 6848 386294 6860
rect 531314 6848 531320 6860
rect 386288 6820 531320 6848
rect 386288 6808 386294 6820
rect 531314 6808 531320 6820
rect 531372 6808 531378 6860
rect 347682 6740 347688 6792
rect 347740 6780 347746 6792
rect 378870 6780 378876 6792
rect 347740 6752 378876 6780
rect 347740 6740 347746 6752
rect 378870 6740 378876 6752
rect 378928 6740 378934 6792
rect 388990 6740 388996 6792
rect 389048 6780 389054 6792
rect 398101 6783 398159 6789
rect 398101 6780 398113 6783
rect 389048 6752 398113 6780
rect 389048 6740 389054 6752
rect 398101 6749 398113 6752
rect 398147 6749 398159 6783
rect 398101 6743 398159 6749
rect 398193 6783 398251 6789
rect 398193 6749 398205 6783
rect 398239 6780 398251 6783
rect 534902 6780 534908 6792
rect 398239 6752 534908 6780
rect 398239 6749 398251 6752
rect 398193 6743 398251 6749
rect 534902 6740 534908 6752
rect 534960 6740 534966 6792
rect 340782 6672 340788 6724
rect 340840 6712 340846 6724
rect 348881 6715 348939 6721
rect 348881 6712 348893 6715
rect 340840 6684 348893 6712
rect 340840 6672 340846 6684
rect 348881 6681 348893 6684
rect 348927 6681 348939 6715
rect 348881 6675 348939 6681
rect 348970 6672 348976 6724
rect 349028 6712 349034 6724
rect 382366 6712 382372 6724
rect 349028 6684 382372 6712
rect 349028 6672 349034 6684
rect 382366 6672 382372 6684
rect 382424 6672 382430 6724
rect 389082 6672 389088 6724
rect 389140 6712 389146 6724
rect 538398 6712 538404 6724
rect 389140 6684 538404 6712
rect 389140 6672 389146 6684
rect 538398 6672 538404 6684
rect 538456 6672 538462 6724
rect 223540 6616 335354 6644
rect 223540 6604 223546 6616
rect 340690 6604 340696 6656
rect 340748 6644 340754 6656
rect 348786 6644 348792 6656
rect 340748 6616 348792 6644
rect 340748 6604 340754 6616
rect 348786 6604 348792 6616
rect 348844 6604 348850 6656
rect 349062 6604 349068 6656
rect 349120 6644 349126 6656
rect 385954 6644 385960 6656
rect 349120 6616 385960 6644
rect 349120 6604 349126 6616
rect 385954 6604 385960 6616
rect 386012 6604 386018 6656
rect 390462 6604 390468 6656
rect 390520 6644 390526 6656
rect 394513 6647 394571 6653
rect 394513 6644 394525 6647
rect 390520 6616 394525 6644
rect 390520 6604 390526 6616
rect 394513 6613 394525 6616
rect 394559 6613 394571 6647
rect 394513 6607 394571 6613
rect 394602 6604 394608 6656
rect 394660 6644 394666 6656
rect 398009 6647 398067 6653
rect 398009 6644 398021 6647
rect 394660 6616 398021 6644
rect 394660 6604 394666 6616
rect 398009 6613 398021 6616
rect 398055 6613 398067 6647
rect 398009 6607 398067 6613
rect 398101 6647 398159 6653
rect 398101 6613 398113 6647
rect 398147 6644 398159 6647
rect 541986 6644 541992 6656
rect 398147 6616 541992 6644
rect 398147 6613 398159 6616
rect 398101 6607 398159 6613
rect 541986 6604 541992 6616
rect 542044 6604 542050 6656
rect 1104 6480 582820 6576
rect 223390 6400 223396 6452
rect 223448 6440 223454 6452
rect 349246 6440 349252 6452
rect 223448 6412 349252 6440
rect 223448 6400 223454 6412
rect 349246 6400 349252 6412
rect 349304 6400 349310 6452
rect 349341 6443 349399 6449
rect 349341 6409 349353 6443
rect 349387 6440 349399 6443
rect 350350 6440 350356 6452
rect 349387 6412 350356 6440
rect 349387 6409 349399 6412
rect 349341 6403 349399 6409
rect 350350 6400 350356 6412
rect 350408 6400 350414 6452
rect 350442 6400 350448 6452
rect 350500 6440 350506 6452
rect 389450 6440 389456 6452
rect 350500 6412 389456 6440
rect 350500 6400 350506 6412
rect 389450 6400 389456 6412
rect 389508 6400 389514 6452
rect 391750 6400 391756 6452
rect 391808 6440 391814 6452
rect 394421 6443 394479 6449
rect 394421 6440 394433 6443
rect 391808 6412 394433 6440
rect 391808 6400 391814 6412
rect 394421 6409 394433 6412
rect 394467 6409 394479 6443
rect 394421 6403 394479 6409
rect 394513 6443 394571 6449
rect 394513 6409 394525 6443
rect 394559 6440 394571 6443
rect 545482 6440 545488 6452
rect 394559 6412 545488 6440
rect 394559 6409 394571 6412
rect 394513 6403 394571 6409
rect 545482 6400 545488 6412
rect 545540 6400 545546 6452
rect 224862 6332 224868 6384
rect 224920 6372 224926 6384
rect 224920 6344 351776 6372
rect 224920 6332 224926 6344
rect 184842 6264 184848 6316
rect 184900 6304 184906 6316
rect 193214 6304 193220 6316
rect 184900 6276 193220 6304
rect 184900 6264 184906 6276
rect 193214 6264 193220 6276
rect 193272 6264 193278 6316
rect 226150 6264 226156 6316
rect 226208 6304 226214 6316
rect 349893 6307 349951 6313
rect 349893 6304 349905 6307
rect 226208 6276 349905 6304
rect 226208 6264 226214 6276
rect 349893 6273 349905 6276
rect 349939 6273 349951 6307
rect 351748 6304 351776 6344
rect 351822 6332 351828 6384
rect 351880 6372 351886 6384
rect 351880 6344 391796 6372
rect 351880 6332 351886 6344
rect 352834 6304 352840 6316
rect 351748 6276 352840 6304
rect 349893 6267 349951 6273
rect 352834 6264 352840 6276
rect 352892 6264 352898 6316
rect 387702 6264 387708 6316
rect 387760 6304 387766 6316
rect 391768 6304 391796 6344
rect 391842 6332 391848 6384
rect 391900 6372 391906 6384
rect 549070 6372 549076 6384
rect 391900 6344 549076 6372
rect 391900 6332 391906 6344
rect 549070 6332 549076 6344
rect 549128 6332 549134 6384
rect 393038 6304 393044 6316
rect 387760 6276 390048 6304
rect 391768 6276 393044 6304
rect 387760 6264 387766 6276
rect 76190 6196 76196 6248
rect 76248 6236 76254 6248
rect 88334 6236 88340 6248
rect 76248 6208 88340 6236
rect 76248 6196 76254 6208
rect 88334 6196 88340 6208
rect 88392 6196 88398 6248
rect 98638 6196 98644 6248
rect 98696 6236 98702 6248
rect 124214 6236 124220 6248
rect 98696 6208 124220 6236
rect 98696 6196 98702 6208
rect 124214 6196 124220 6208
rect 124272 6196 124278 6248
rect 188982 6196 188988 6248
rect 189040 6236 189046 6248
rect 210970 6236 210976 6248
rect 189040 6208 210976 6236
rect 189040 6196 189046 6208
rect 210970 6196 210976 6208
rect 211028 6196 211034 6248
rect 226242 6196 226248 6248
rect 226300 6236 226306 6248
rect 359918 6236 359924 6248
rect 226300 6208 359924 6236
rect 226300 6196 226306 6208
rect 359918 6196 359924 6208
rect 359976 6196 359982 6248
rect 380802 6196 380808 6248
rect 380860 6236 380866 6248
rect 388441 6239 388499 6245
rect 388441 6236 388453 6239
rect 380860 6208 388453 6236
rect 380860 6196 380866 6208
rect 388441 6205 388453 6208
rect 388487 6205 388499 6239
rect 390020 6236 390048 6276
rect 393038 6264 393044 6276
rect 393096 6264 393102 6316
rect 393222 6264 393228 6316
rect 393280 6304 393286 6316
rect 394789 6307 394847 6313
rect 393280 6276 394740 6304
rect 393280 6264 393286 6276
rect 394602 6236 394608 6248
rect 390020 6208 394608 6236
rect 388441 6199 388499 6205
rect 394602 6196 394608 6208
rect 394660 6196 394666 6248
rect 394712 6236 394740 6276
rect 394789 6273 394801 6307
rect 394835 6304 394847 6307
rect 552658 6304 552664 6316
rect 394835 6276 552664 6304
rect 394835 6273 394847 6276
rect 394789 6267 394847 6273
rect 552658 6264 552664 6276
rect 552716 6264 552722 6316
rect 463697 6239 463755 6245
rect 463697 6236 463709 6239
rect 394712 6208 463709 6236
rect 463697 6205 463709 6208
rect 463743 6205 463755 6239
rect 463878 6236 463884 6248
rect 463839 6208 463884 6236
rect 463697 6199 463755 6205
rect 463878 6196 463884 6208
rect 463936 6196 463942 6248
rect 463973 6239 464031 6245
rect 463973 6205 463985 6239
rect 464019 6236 464031 6239
rect 556154 6236 556160 6248
rect 464019 6208 556160 6236
rect 464019 6205 464031 6208
rect 463973 6199 464031 6205
rect 556154 6196 556160 6208
rect 556212 6196 556218 6248
rect 26510 6128 26516 6180
rect 26568 6168 26574 6180
rect 75914 6168 75920 6180
rect 26568 6140 75920 6168
rect 26568 6128 26574 6140
rect 75914 6128 75920 6140
rect 75972 6128 75978 6180
rect 77386 6128 77392 6180
rect 77444 6168 77450 6180
rect 118694 6168 118700 6180
rect 77444 6140 118700 6168
rect 77444 6128 77450 6140
rect 118694 6128 118700 6140
rect 118752 6128 118758 6180
rect 125870 6128 125876 6180
rect 125928 6168 125934 6180
rect 165614 6168 165620 6180
rect 125928 6140 165620 6168
rect 125928 6128 125934 6140
rect 165614 6128 165620 6140
rect 165672 6128 165678 6180
rect 191650 6128 191656 6180
rect 191708 6168 191714 6180
rect 221550 6168 221556 6180
rect 191708 6140 221556 6168
rect 191708 6128 191714 6140
rect 221550 6128 221556 6140
rect 221608 6128 221614 6180
rect 227622 6128 227628 6180
rect 227680 6168 227686 6180
rect 363506 6168 363512 6180
rect 227680 6140 363512 6168
rect 227680 6128 227686 6140
rect 363506 6128 363512 6140
rect 363564 6128 363570 6180
rect 379422 6128 379428 6180
rect 379480 6168 379486 6180
rect 502150 6168 502156 6180
rect 379480 6140 502156 6168
rect 379480 6128 379486 6140
rect 502150 6128 502156 6140
rect 502208 6128 502214 6180
rect 502245 6171 502303 6177
rect 502245 6137 502257 6171
rect 502291 6168 502303 6171
rect 559742 6168 559748 6180
rect 502291 6140 559748 6168
rect 502291 6137 502303 6140
rect 502245 6131 502303 6137
rect 559742 6128 559748 6140
rect 559800 6128 559806 6180
rect 297266 6060 297272 6112
rect 297324 6100 297330 6112
rect 325694 6100 325700 6112
rect 297324 6072 325700 6100
rect 297324 6060 297330 6072
rect 325694 6060 325700 6072
rect 325752 6060 325758 6112
rect 346302 6060 346308 6112
rect 346360 6100 346366 6112
rect 371694 6100 371700 6112
rect 346360 6072 371700 6100
rect 346360 6060 346366 6072
rect 371694 6060 371700 6072
rect 371752 6060 371758 6112
rect 386138 6060 386144 6112
rect 386196 6100 386202 6112
rect 527818 6100 527824 6112
rect 386196 6072 527824 6100
rect 386196 6060 386202 6072
rect 527818 6060 527824 6072
rect 527876 6060 527882 6112
rect 1104 5936 582820 6032
rect 300762 5856 300768 5908
rect 300820 5896 300826 5908
rect 327074 5896 327080 5908
rect 300820 5868 327080 5896
rect 300820 5856 300826 5868
rect 327074 5856 327080 5868
rect 327132 5856 327138 5908
rect 344922 5856 344928 5908
rect 344980 5896 344986 5908
rect 368198 5896 368204 5908
rect 344980 5868 368204 5896
rect 344980 5856 344986 5868
rect 368198 5856 368204 5868
rect 368256 5856 368262 5908
rect 384942 5856 384948 5908
rect 385000 5896 385006 5908
rect 524230 5896 524236 5908
rect 385000 5868 524236 5896
rect 385000 5856 385006 5868
rect 524230 5856 524236 5868
rect 524288 5856 524294 5908
rect 304350 5788 304356 5840
rect 304408 5828 304414 5840
rect 327166 5828 327172 5840
rect 304408 5800 327172 5828
rect 304408 5788 304414 5800
rect 327166 5788 327172 5800
rect 327224 5788 327230 5840
rect 327721 5831 327779 5837
rect 327721 5797 327733 5831
rect 327767 5828 327779 5831
rect 331214 5828 331220 5840
rect 327767 5800 331220 5828
rect 327767 5797 327779 5800
rect 327721 5791 327779 5797
rect 331214 5788 331220 5800
rect 331272 5788 331278 5840
rect 337930 5788 337936 5840
rect 337988 5828 337994 5840
rect 343358 5828 343364 5840
rect 337988 5800 343364 5828
rect 337988 5788 337994 5800
rect 343358 5788 343364 5800
rect 343416 5788 343422 5840
rect 343542 5788 343548 5840
rect 343600 5828 343606 5840
rect 364610 5828 364616 5840
rect 343600 5800 364616 5828
rect 343600 5788 343606 5800
rect 364610 5788 364616 5800
rect 364668 5788 364674 5840
rect 383562 5788 383568 5840
rect 383620 5828 383626 5840
rect 520734 5828 520740 5840
rect 383620 5800 520740 5828
rect 383620 5788 383626 5800
rect 520734 5788 520740 5800
rect 520792 5788 520798 5840
rect 520918 5788 520924 5840
rect 520976 5828 520982 5840
rect 580166 5828 580172 5840
rect 520976 5800 580172 5828
rect 520976 5788 520982 5800
rect 580166 5788 580172 5800
rect 580224 5788 580230 5840
rect 307938 5720 307944 5772
rect 307996 5760 308002 5772
rect 328454 5760 328460 5772
rect 307996 5732 328460 5760
rect 307996 5720 308002 5732
rect 328454 5720 328460 5732
rect 328512 5720 328518 5772
rect 339402 5720 339408 5772
rect 339460 5760 339466 5772
rect 339460 5732 343404 5760
rect 339460 5720 339466 5732
rect 315022 5652 315028 5704
rect 315080 5692 315086 5704
rect 320729 5695 320787 5701
rect 320729 5692 320741 5695
rect 315080 5664 320741 5692
rect 315080 5652 315086 5664
rect 320729 5661 320741 5664
rect 320775 5661 320787 5695
rect 329834 5692 329840 5704
rect 320729 5655 320787 5661
rect 320836 5664 329840 5692
rect 209409 5627 209467 5633
rect 209409 5593 209421 5627
rect 209455 5624 209467 5627
rect 219621 5627 219679 5633
rect 219621 5624 219633 5627
rect 209455 5596 219633 5624
rect 209455 5593 209467 5596
rect 209409 5587 209467 5593
rect 219621 5593 219633 5596
rect 219667 5593 219679 5627
rect 219621 5587 219679 5593
rect 277029 5627 277087 5633
rect 277029 5593 277041 5627
rect 277075 5624 277087 5627
rect 282822 5624 282828 5636
rect 277075 5596 282828 5624
rect 277075 5593 277087 5596
rect 277029 5587 277087 5593
rect 282822 5584 282828 5596
rect 282880 5584 282886 5636
rect 311434 5584 311440 5636
rect 311492 5624 311498 5636
rect 320836 5624 320864 5664
rect 329834 5652 329840 5664
rect 329892 5652 329898 5704
rect 343376 5692 343404 5732
rect 343450 5720 343456 5772
rect 343508 5760 343514 5772
rect 361114 5760 361120 5772
rect 343508 5732 361120 5760
rect 343508 5720 343514 5732
rect 361114 5720 361120 5732
rect 361172 5720 361178 5772
rect 383470 5720 383476 5772
rect 383528 5760 383534 5772
rect 517146 5760 517152 5772
rect 383528 5732 517152 5760
rect 383528 5720 383534 5732
rect 517146 5720 517152 5732
rect 517204 5720 517210 5772
rect 346946 5692 346952 5704
rect 343376 5664 346952 5692
rect 346946 5652 346952 5664
rect 347004 5652 347010 5704
rect 357526 5692 357532 5704
rect 349816 5664 357532 5692
rect 311492 5596 320864 5624
rect 320928 5596 327856 5624
rect 311492 5584 311498 5596
rect 86862 5516 86868 5568
rect 86920 5556 86926 5568
rect 91094 5556 91100 5568
rect 86920 5528 91100 5556
rect 86920 5516 86926 5528
rect 91094 5516 91100 5528
rect 91152 5516 91158 5568
rect 184198 5516 184204 5568
rect 184256 5556 184262 5568
rect 189718 5556 189724 5568
rect 184256 5528 189724 5556
rect 184256 5516 184262 5528
rect 189718 5516 189724 5528
rect 189776 5516 189782 5568
rect 209501 5559 209559 5565
rect 209501 5525 209513 5559
rect 209547 5556 209559 5559
rect 219713 5559 219771 5565
rect 219713 5556 219725 5559
rect 209547 5528 219725 5556
rect 209547 5525 209559 5528
rect 209501 5519 209559 5525
rect 219713 5525 219725 5528
rect 219759 5525 219771 5559
rect 219713 5519 219771 5525
rect 275922 5516 275928 5568
rect 275980 5556 275986 5568
rect 279697 5559 279755 5565
rect 279697 5556 279709 5559
rect 275980 5528 279709 5556
rect 275980 5516 275986 5528
rect 279697 5525 279709 5528
rect 279743 5525 279755 5559
rect 279697 5519 279755 5525
rect 282641 5559 282699 5565
rect 282641 5525 282653 5559
rect 282687 5556 282699 5559
rect 316034 5556 316040 5568
rect 282687 5528 316040 5556
rect 282687 5525 282699 5528
rect 282641 5519 282699 5525
rect 316034 5516 316040 5528
rect 316092 5516 316098 5568
rect 318518 5516 318524 5568
rect 318576 5556 318582 5568
rect 320637 5559 320695 5565
rect 320637 5556 320649 5559
rect 318576 5528 320649 5556
rect 318576 5516 318582 5528
rect 320637 5525 320649 5528
rect 320683 5525 320695 5559
rect 320637 5519 320695 5525
rect 320729 5559 320787 5565
rect 320729 5525 320741 5559
rect 320775 5556 320787 5559
rect 320928 5556 320956 5596
rect 320775 5528 320956 5556
rect 321005 5559 321063 5565
rect 320775 5525 320787 5528
rect 320729 5519 320787 5525
rect 321005 5525 321017 5559
rect 321051 5556 321063 5559
rect 327721 5559 327779 5565
rect 327721 5556 327733 5559
rect 321051 5528 327733 5556
rect 321051 5525 321063 5528
rect 321005 5519 321063 5525
rect 327721 5525 327733 5528
rect 327767 5525 327779 5559
rect 327828 5556 327856 5596
rect 329190 5584 329196 5636
rect 329248 5624 329254 5636
rect 334066 5624 334072 5636
rect 329248 5596 334072 5624
rect 329248 5584 329254 5596
rect 334066 5584 334072 5596
rect 334124 5584 334130 5636
rect 334158 5584 334164 5636
rect 334216 5624 334222 5636
rect 334216 5596 335354 5624
rect 334216 5584 334222 5596
rect 329926 5556 329932 5568
rect 327828 5528 329932 5556
rect 327721 5519 327779 5525
rect 329926 5516 329932 5528
rect 329984 5516 329990 5568
rect 332686 5516 332692 5568
rect 332744 5556 332750 5568
rect 333974 5556 333980 5568
rect 332744 5528 333980 5556
rect 332744 5516 332750 5528
rect 333974 5516 333980 5528
rect 334032 5516 334038 5568
rect 335326 5556 335354 5596
rect 338022 5584 338028 5636
rect 338080 5624 338086 5636
rect 339862 5624 339868 5636
rect 338080 5596 339868 5624
rect 338080 5584 338086 5596
rect 339862 5584 339868 5596
rect 339920 5584 339926 5636
rect 342162 5584 342168 5636
rect 342220 5624 342226 5636
rect 349816 5624 349844 5664
rect 357526 5652 357532 5664
rect 357584 5652 357590 5704
rect 382182 5652 382188 5704
rect 382240 5692 382246 5704
rect 513558 5692 513564 5704
rect 382240 5664 513564 5692
rect 382240 5652 382246 5664
rect 513558 5652 513564 5664
rect 513616 5652 513622 5704
rect 342220 5596 349844 5624
rect 349893 5627 349951 5633
rect 342220 5584 342226 5596
rect 349893 5593 349905 5627
rect 349939 5624 349951 5627
rect 356330 5624 356336 5636
rect 349939 5596 356336 5624
rect 349939 5593 349951 5596
rect 349893 5587 349951 5593
rect 356330 5584 356336 5596
rect 356388 5584 356394 5636
rect 380710 5584 380716 5636
rect 380768 5624 380774 5636
rect 510062 5624 510068 5636
rect 380768 5596 510068 5624
rect 380768 5584 380774 5596
rect 510062 5584 510068 5596
rect 510120 5584 510126 5636
rect 383654 5556 383660 5568
rect 335326 5528 383660 5556
rect 383654 5516 383660 5528
rect 383712 5516 383718 5568
rect 388441 5559 388499 5565
rect 388441 5525 388453 5559
rect 388487 5556 388499 5559
rect 499666 5556 499672 5568
rect 388487 5528 499672 5556
rect 388487 5525 388499 5528
rect 388441 5519 388499 5525
rect 499666 5516 499672 5528
rect 499724 5516 499730 5568
rect 499758 5516 499764 5568
rect 499816 5556 499822 5568
rect 509329 5559 509387 5565
rect 509329 5556 509341 5559
rect 499816 5528 509341 5556
rect 499816 5516 499822 5528
rect 509329 5525 509341 5528
rect 509375 5525 509387 5559
rect 509329 5519 509387 5525
rect 514570 5516 514576 5568
rect 514628 5556 514634 5568
rect 521933 5559 521991 5565
rect 521933 5556 521945 5559
rect 514628 5528 521945 5556
rect 514628 5516 514634 5528
rect 521933 5525 521945 5528
rect 521979 5525 521991 5559
rect 521933 5519 521991 5525
rect 1104 5392 582820 5488
rect 63218 5312 63224 5364
rect 63276 5352 63282 5364
rect 114554 5352 114560 5364
rect 63276 5324 114560 5352
rect 63276 5312 63282 5324
rect 114554 5312 114560 5324
rect 114612 5312 114618 5364
rect 200022 5312 200028 5364
rect 200080 5352 200086 5364
rect 257062 5352 257068 5364
rect 200080 5324 257068 5352
rect 200080 5312 200086 5324
rect 257062 5312 257068 5324
rect 257120 5312 257126 5364
rect 274450 5312 274456 5364
rect 274508 5352 274514 5364
rect 277029 5355 277087 5361
rect 277029 5352 277041 5355
rect 274508 5324 277041 5352
rect 274508 5312 274514 5324
rect 277029 5321 277041 5324
rect 277075 5321 277087 5355
rect 277029 5315 277087 5321
rect 277118 5312 277124 5364
rect 277176 5352 277182 5364
rect 277176 5324 278360 5352
rect 277176 5312 277182 5324
rect 56042 5244 56048 5296
rect 56100 5284 56106 5296
rect 113266 5284 113272 5296
rect 56100 5256 113272 5284
rect 56100 5244 56106 5256
rect 113266 5244 113272 5256
rect 113324 5244 113330 5296
rect 201402 5244 201408 5296
rect 201460 5284 201466 5296
rect 205266 5284 205272 5296
rect 201460 5256 205272 5284
rect 201460 5244 201466 5256
rect 205266 5244 205272 5256
rect 205324 5244 205330 5296
rect 205542 5244 205548 5296
rect 205600 5284 205606 5296
rect 209409 5287 209467 5293
rect 209409 5284 209421 5287
rect 205600 5256 209421 5284
rect 205600 5244 205606 5256
rect 209409 5253 209421 5256
rect 209455 5253 209467 5287
rect 209409 5247 209467 5253
rect 209593 5287 209651 5293
rect 209593 5253 209605 5287
rect 209639 5284 209651 5287
rect 267734 5284 267740 5296
rect 209639 5256 267740 5284
rect 209639 5253 209651 5256
rect 209593 5247 209651 5253
rect 267734 5244 267740 5256
rect 267792 5244 267798 5296
rect 274542 5244 274548 5296
rect 274600 5284 274606 5296
rect 278225 5287 278283 5293
rect 278225 5284 278237 5287
rect 274600 5256 278237 5284
rect 274600 5244 274606 5256
rect 278225 5253 278237 5256
rect 278271 5253 278283 5287
rect 278225 5247 278283 5253
rect 48958 5176 48964 5228
rect 49016 5216 49022 5228
rect 110414 5216 110420 5228
rect 49016 5188 110420 5216
rect 49016 5176 49022 5188
rect 110414 5176 110420 5188
rect 110472 5176 110478 5228
rect 202782 5176 202788 5228
rect 202840 5216 202846 5228
rect 205358 5216 205364 5228
rect 202840 5188 205364 5216
rect 202840 5176 202846 5188
rect 205358 5176 205364 5188
rect 205416 5176 205422 5228
rect 205450 5176 205456 5228
rect 205508 5216 205514 5228
rect 209501 5219 209559 5225
rect 209501 5216 209513 5219
rect 205508 5188 209513 5216
rect 205508 5176 205514 5188
rect 209501 5185 209513 5188
rect 209547 5185 209559 5219
rect 209501 5179 209559 5185
rect 209685 5219 209743 5225
rect 209685 5185 209697 5219
rect 209731 5216 209743 5219
rect 271230 5216 271236 5228
rect 209731 5188 271236 5216
rect 209731 5185 209743 5188
rect 209685 5179 209743 5185
rect 271230 5176 271236 5188
rect 271288 5176 271294 5228
rect 271782 5176 271788 5228
rect 271840 5216 271846 5228
rect 278133 5219 278191 5225
rect 278133 5216 278145 5219
rect 271840 5188 278145 5216
rect 271840 5176 271846 5188
rect 278133 5185 278145 5188
rect 278179 5185 278191 5219
rect 278332 5216 278360 5324
rect 278682 5312 278688 5364
rect 278740 5352 278746 5364
rect 282641 5355 282699 5361
rect 282641 5352 282653 5355
rect 278740 5324 282653 5352
rect 278740 5312 278746 5324
rect 282641 5321 282653 5324
rect 282687 5321 282699 5355
rect 544378 5352 544384 5364
rect 282641 5315 282699 5321
rect 282748 5324 544384 5352
rect 278409 5287 278467 5293
rect 278409 5253 278421 5287
rect 278455 5284 278467 5287
rect 282748 5284 282776 5324
rect 544378 5312 544384 5324
rect 544436 5312 544442 5364
rect 278455 5256 282776 5284
rect 278455 5253 278467 5256
rect 278409 5247 278467 5253
rect 282822 5244 282828 5296
rect 282880 5284 282886 5296
rect 547874 5284 547880 5296
rect 282880 5256 547880 5284
rect 282880 5244 282886 5256
rect 547874 5244 547880 5256
rect 547932 5244 547938 5296
rect 279697 5219 279755 5225
rect 278332 5188 279648 5216
rect 278133 5179 278191 5185
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 70394 5148 70400 5160
rect 1728 5120 70400 5148
rect 1728 5108 1734 5120
rect 70394 5108 70400 5120
rect 70452 5108 70458 5160
rect 97902 5108 97908 5160
rect 97960 5148 97966 5160
rect 108114 5148 108120 5160
rect 97960 5120 108120 5148
rect 97960 5108 97966 5120
rect 108114 5108 108120 5120
rect 108172 5108 108178 5160
rect 191742 5108 191748 5160
rect 191800 5148 191806 5160
rect 219434 5148 219440 5160
rect 191800 5120 219440 5148
rect 191800 5108 191806 5120
rect 219434 5108 219440 5120
rect 219492 5108 219498 5160
rect 219713 5151 219771 5157
rect 219713 5117 219725 5151
rect 219759 5148 219771 5151
rect 274818 5148 274824 5160
rect 219759 5120 274824 5148
rect 219759 5117 219771 5120
rect 219713 5111 219771 5117
rect 274818 5108 274824 5120
rect 274876 5108 274882 5160
rect 277210 5108 277216 5160
rect 277268 5148 277274 5160
rect 279620 5148 279648 5188
rect 279697 5185 279709 5219
rect 279743 5216 279755 5219
rect 551462 5216 551468 5228
rect 279743 5188 551468 5216
rect 279743 5185 279755 5188
rect 279697 5179 279755 5185
rect 551462 5176 551468 5188
rect 551520 5176 551526 5228
rect 554958 5148 554964 5160
rect 277268 5120 279556 5148
rect 279620 5120 554964 5148
rect 277268 5108 277274 5120
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 71774 5080 71780 5092
rect 2924 5052 71780 5080
rect 2924 5040 2930 5052
rect 71774 5040 71780 5052
rect 71832 5040 71838 5092
rect 99190 5040 99196 5092
rect 99248 5080 99254 5092
rect 115198 5080 115204 5092
rect 99248 5052 115204 5080
rect 99248 5040 99254 5052
rect 115198 5040 115204 5052
rect 115256 5040 115262 5092
rect 193122 5040 193128 5092
rect 193180 5080 193186 5092
rect 219529 5083 219587 5089
rect 219529 5080 219541 5083
rect 193180 5052 219541 5080
rect 193180 5040 193186 5052
rect 219529 5049 219541 5052
rect 219575 5049 219587 5083
rect 219529 5043 219587 5049
rect 219621 5083 219679 5089
rect 219621 5049 219633 5083
rect 219667 5080 219679 5083
rect 278314 5080 278320 5092
rect 219667 5052 278320 5080
rect 219667 5049 219679 5052
rect 219621 5043 219679 5049
rect 278314 5040 278320 5052
rect 278372 5040 278378 5092
rect 279528 5080 279556 5120
rect 554958 5108 554964 5120
rect 555016 5108 555022 5160
rect 558546 5080 558552 5092
rect 279528 5052 558552 5080
rect 558546 5040 558552 5052
rect 558604 5040 558610 5092
rect 566 4972 572 5024
rect 624 5012 630 5024
rect 70486 5012 70492 5024
rect 624 4984 70492 5012
rect 624 4972 630 4984
rect 70486 4972 70492 4984
rect 70544 4972 70550 5024
rect 100662 4972 100668 5024
rect 100720 5012 100726 5024
rect 118786 5012 118792 5024
rect 100720 4984 118792 5012
rect 100720 4972 100726 4984
rect 118786 4972 118792 4984
rect 118844 4972 118850 5024
rect 204162 4972 204168 5024
rect 204220 5012 204226 5024
rect 209501 5015 209559 5021
rect 209501 5012 209513 5015
rect 204220 4984 209513 5012
rect 204220 4972 204226 4984
rect 209501 4981 209513 4984
rect 209547 4981 209559 5015
rect 209501 4975 209559 4981
rect 209682 4972 209688 5024
rect 209740 5012 209746 5024
rect 260650 5012 260656 5024
rect 209740 4984 260656 5012
rect 209740 4972 209746 4984
rect 260650 4972 260656 4984
rect 260708 4972 260714 5024
rect 266262 4972 266268 5024
rect 266320 5012 266326 5024
rect 509234 5012 509240 5024
rect 266320 4984 509240 5012
rect 266320 4972 266326 4984
rect 509234 4972 509240 4984
rect 509292 4972 509298 5024
rect 509329 5015 509387 5021
rect 509329 4981 509341 5015
rect 509375 5012 509387 5015
rect 562042 5012 562048 5024
rect 509375 4984 562048 5012
rect 509375 4981 509387 4984
rect 509329 4975 509387 4981
rect 562042 4972 562048 4984
rect 562100 4972 562106 5024
rect 1104 4848 582820 4944
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 100754 4808 100760 4820
rect 4120 4780 100760 4808
rect 4120 4768 4126 4780
rect 100754 4768 100760 4780
rect 100812 4768 100818 4820
rect 102042 4768 102048 4820
rect 102100 4808 102106 4820
rect 122282 4808 122288 4820
rect 102100 4780 122288 4808
rect 102100 4768 102106 4780
rect 122282 4768 122288 4780
rect 122340 4768 122346 4820
rect 202690 4768 202696 4820
rect 202748 4808 202754 4820
rect 209409 4811 209467 4817
rect 209409 4808 209421 4811
rect 202748 4780 209421 4808
rect 202748 4768 202754 4780
rect 209409 4777 209421 4780
rect 209455 4777 209467 4811
rect 209409 4771 209467 4777
rect 209590 4768 209596 4820
rect 209648 4808 209654 4820
rect 264146 4808 264152 4820
rect 209648 4780 264152 4808
rect 209648 4768 209654 4780
rect 264146 4768 264152 4780
rect 264204 4768 264210 4820
rect 266170 4768 266176 4820
rect 266228 4808 266234 4820
rect 480254 4808 480260 4820
rect 266228 4780 480260 4808
rect 266228 4768 266234 4780
rect 480254 4768 480260 4780
rect 480312 4768 480318 4820
rect 480346 4768 480352 4820
rect 480404 4808 480410 4820
rect 489822 4808 489828 4820
rect 480404 4780 489828 4808
rect 480404 4768 480410 4780
rect 489822 4768 489828 4780
rect 489880 4768 489886 4820
rect 489914 4768 489920 4820
rect 489972 4808 489978 4820
rect 499390 4808 499396 4820
rect 489972 4780 499396 4808
rect 489972 4768 489978 4780
rect 499390 4768 499396 4780
rect 499448 4768 499454 4820
rect 499482 4768 499488 4820
rect 499540 4808 499546 4820
rect 509237 4811 509295 4817
rect 509237 4808 509249 4811
rect 499540 4780 509249 4808
rect 499540 4768 499546 4780
rect 509237 4777 509249 4780
rect 509283 4777 509295 4811
rect 509237 4771 509295 4777
rect 509329 4811 509387 4817
rect 509329 4777 509341 4811
rect 509375 4808 509387 4811
rect 565630 4808 565636 4820
rect 509375 4780 565636 4808
rect 509375 4777 509387 4780
rect 509329 4771 509387 4777
rect 565630 4768 565636 4780
rect 565688 4768 565694 4820
rect 47854 4700 47860 4752
rect 47912 4740 47918 4752
rect 81434 4740 81440 4752
rect 47912 4712 81440 4740
rect 47912 4700 47918 4712
rect 81434 4700 81440 4712
rect 81492 4700 81498 4752
rect 99282 4700 99288 4752
rect 99340 4740 99346 4752
rect 111610 4740 111616 4752
rect 99340 4712 111616 4740
rect 99340 4700 99346 4712
rect 111610 4700 111616 4712
rect 111668 4700 111674 4752
rect 199930 4700 199936 4752
rect 199988 4740 199994 4752
rect 253474 4740 253480 4752
rect 199988 4712 253480 4740
rect 199988 4700 199994 4712
rect 253474 4700 253480 4712
rect 253532 4700 253538 4752
rect 271690 4700 271696 4752
rect 271748 4740 271754 4752
rect 277857 4743 277915 4749
rect 277857 4740 277869 4743
rect 271748 4712 277869 4740
rect 271748 4700 271754 4712
rect 277857 4709 277869 4712
rect 277903 4709 277915 4743
rect 540790 4740 540796 4752
rect 277857 4703 277915 4709
rect 277964 4712 540796 4740
rect 51350 4632 51356 4684
rect 51408 4672 51414 4684
rect 81526 4672 81532 4684
rect 51408 4644 81532 4672
rect 51408 4632 51414 4644
rect 81526 4632 81532 4644
rect 81584 4632 81590 4684
rect 96154 4632 96160 4684
rect 96212 4672 96218 4684
rect 104526 4672 104532 4684
rect 96212 4644 104532 4672
rect 96212 4632 96218 4644
rect 104526 4632 104532 4644
rect 104584 4632 104590 4684
rect 198642 4632 198648 4684
rect 198700 4672 198706 4684
rect 249978 4672 249984 4684
rect 198700 4644 249984 4672
rect 198700 4632 198706 4644
rect 249978 4632 249984 4644
rect 250036 4632 250042 4684
rect 54938 4564 54944 4616
rect 54996 4604 55002 4616
rect 82814 4604 82820 4616
rect 54996 4576 82820 4604
rect 54996 4564 55002 4576
rect 82814 4564 82820 4576
rect 82872 4564 82878 4616
rect 197262 4564 197268 4616
rect 197320 4604 197326 4616
rect 246390 4604 246396 4616
rect 197320 4576 246396 4604
rect 197320 4564 197326 4576
rect 246390 4564 246396 4576
rect 246448 4564 246454 4616
rect 273162 4564 273168 4616
rect 273220 4604 273226 4616
rect 277964 4604 277992 4712
rect 540790 4700 540796 4712
rect 540848 4700 540854 4752
rect 278041 4675 278099 4681
rect 278041 4641 278053 4675
rect 278087 4672 278099 4675
rect 537202 4672 537208 4684
rect 278087 4644 537208 4672
rect 278087 4641 278099 4644
rect 278041 4635 278099 4641
rect 537202 4632 537208 4644
rect 537260 4632 537266 4684
rect 273220 4576 277992 4604
rect 278133 4607 278191 4613
rect 273220 4564 273226 4576
rect 278133 4573 278145 4607
rect 278179 4604 278191 4607
rect 533706 4604 533712 4616
rect 278179 4576 533712 4604
rect 278179 4573 278191 4576
rect 278133 4567 278191 4573
rect 533706 4564 533712 4576
rect 533764 4564 533770 4616
rect 65518 4496 65524 4548
rect 65576 4536 65582 4548
rect 85574 4536 85580 4548
rect 65576 4508 85580 4536
rect 65576 4496 65582 4508
rect 85574 4496 85580 4508
rect 85632 4496 85638 4548
rect 197170 4496 197176 4548
rect 197228 4536 197234 4548
rect 242894 4536 242900 4548
rect 197228 4508 242900 4536
rect 197228 4496 197234 4508
rect 242894 4496 242900 4508
rect 242952 4496 242958 4548
rect 270402 4496 270408 4548
rect 270460 4536 270466 4548
rect 530118 4536 530124 4548
rect 270460 4508 530124 4536
rect 270460 4496 270466 4508
rect 530118 4496 530124 4508
rect 530176 4496 530182 4548
rect 69106 4428 69112 4480
rect 69164 4468 69170 4480
rect 86954 4468 86960 4480
rect 69164 4440 86960 4468
rect 69164 4428 69170 4440
rect 86954 4428 86960 4440
rect 87012 4428 87018 4480
rect 195882 4428 195888 4480
rect 195940 4468 195946 4480
rect 239306 4468 239312 4480
rect 195940 4440 239312 4468
rect 195940 4428 195946 4440
rect 239306 4428 239312 4440
rect 239364 4428 239370 4480
rect 268930 4428 268936 4480
rect 268988 4468 268994 4480
rect 526622 4468 526628 4480
rect 268988 4440 526628 4468
rect 268988 4428 268994 4440
rect 526622 4428 526628 4440
rect 526680 4428 526686 4480
rect 1104 4304 582820 4400
rect 96430 4224 96436 4276
rect 96488 4264 96494 4276
rect 101030 4264 101036 4276
rect 96488 4236 101036 4264
rect 96488 4224 96494 4236
rect 101030 4224 101036 4236
rect 101088 4224 101094 4276
rect 194226 4224 194232 4276
rect 194284 4264 194290 4276
rect 235718 4264 235724 4276
rect 194284 4236 235724 4264
rect 194284 4224 194290 4236
rect 235718 4224 235724 4236
rect 235776 4224 235782 4276
rect 269022 4224 269028 4276
rect 269080 4264 269086 4276
rect 523034 4264 523040 4276
rect 269080 4236 523040 4264
rect 269080 4224 269086 4236
rect 523034 4224 523040 4236
rect 523092 4224 523098 4276
rect 95142 4156 95148 4208
rect 95200 4196 95206 4208
rect 97442 4196 97448 4208
rect 95200 4168 97448 4196
rect 95200 4156 95206 4168
rect 97442 4156 97448 4168
rect 97500 4156 97506 4208
rect 123205 4199 123263 4205
rect 123205 4165 123217 4199
rect 123251 4196 123263 4199
rect 128541 4199 128599 4205
rect 128541 4196 128553 4199
rect 123251 4168 128553 4196
rect 123251 4165 123263 4168
rect 123205 4159 123263 4165
rect 128541 4165 128553 4168
rect 128587 4165 128599 4199
rect 128541 4159 128599 4165
rect 132773 4199 132831 4205
rect 132773 4165 132785 4199
rect 132819 4196 132831 4199
rect 135346 4196 135352 4208
rect 132819 4168 135352 4196
rect 132819 4165 132831 4168
rect 132773 4159 132831 4165
rect 135346 4156 135352 4168
rect 135404 4156 135410 4208
rect 194318 4156 194324 4208
rect 194376 4196 194382 4208
rect 232222 4196 232228 4208
rect 194376 4168 232228 4196
rect 194376 4156 194382 4168
rect 232222 4156 232228 4168
rect 232280 4156 232286 4208
rect 267642 4156 267648 4208
rect 267700 4196 267706 4208
rect 519538 4196 519544 4208
rect 267700 4168 519544 4196
rect 267700 4156 267706 4168
rect 519538 4156 519544 4168
rect 519596 4156 519602 4208
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7558 4128 7564 4140
rect 6512 4100 7564 4128
rect 6512 4088 6518 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 149054 4128 149060 4140
rect 85724 4100 149060 4128
rect 85724 4088 85730 4100
rect 149054 4088 149060 4100
rect 149112 4088 149118 4140
rect 158898 4088 158904 4140
rect 158956 4128 158962 4140
rect 160002 4128 160008 4140
rect 158956 4100 160008 4128
rect 158956 4088 158962 4100
rect 160002 4088 160008 4100
rect 160060 4088 160066 4140
rect 164878 4088 164884 4140
rect 164936 4128 164942 4140
rect 165522 4128 165528 4140
rect 164936 4100 165528 4128
rect 164936 4088 164942 4100
rect 165522 4088 165528 4100
rect 165580 4088 165586 4140
rect 219529 4131 219587 4137
rect 219529 4097 219541 4131
rect 219575 4128 219587 4131
rect 228726 4128 228732 4140
rect 219575 4100 228732 4128
rect 219575 4097 219587 4100
rect 219529 4091 219587 4097
rect 228726 4088 228732 4100
rect 228784 4088 228790 4140
rect 273622 4088 273628 4140
rect 273680 4128 273686 4140
rect 274358 4128 274364 4140
rect 273680 4100 274364 4128
rect 273680 4088 273686 4100
rect 274358 4088 274364 4100
rect 274416 4088 274422 4140
rect 277210 4088 277216 4140
rect 277268 4128 277274 4140
rect 278038 4128 278044 4140
rect 277268 4100 278044 4128
rect 277268 4088 277274 4100
rect 278038 4088 278044 4100
rect 278096 4088 278102 4140
rect 283098 4088 283104 4140
rect 283156 4128 283162 4140
rect 284202 4128 284208 4140
rect 283156 4100 284208 4128
rect 283156 4088 283162 4100
rect 284202 4088 284208 4100
rect 284260 4088 284266 4140
rect 284294 4088 284300 4140
rect 284352 4128 284358 4140
rect 285582 4128 285588 4140
rect 284352 4100 285588 4128
rect 284352 4088 284358 4100
rect 285582 4088 285588 4100
rect 285640 4088 285646 4140
rect 287790 4088 287796 4140
rect 287848 4128 287854 4140
rect 288342 4128 288348 4140
rect 287848 4100 288348 4128
rect 287848 4088 287854 4100
rect 288342 4088 288348 4100
rect 288400 4088 288406 4140
rect 291378 4088 291384 4140
rect 291436 4128 291442 4140
rect 292482 4128 292488 4140
rect 291436 4100 292488 4128
rect 291436 4088 291442 4100
rect 292482 4088 292488 4100
rect 292540 4088 292546 4140
rect 298462 4088 298468 4140
rect 298520 4128 298526 4140
rect 299382 4128 299388 4140
rect 298520 4100 299388 4128
rect 298520 4088 298526 4100
rect 299382 4088 299388 4100
rect 299440 4088 299446 4140
rect 305546 4088 305552 4140
rect 305604 4128 305610 4140
rect 308490 4128 308496 4140
rect 305604 4100 308496 4128
rect 305604 4088 305610 4100
rect 308490 4088 308496 4100
rect 308548 4088 308554 4140
rect 309042 4088 309048 4140
rect 309100 4128 309106 4140
rect 309778 4128 309784 4140
rect 309100 4100 309784 4128
rect 309100 4088 309106 4100
rect 309778 4088 309784 4100
rect 309836 4088 309842 4140
rect 383654 4128 383660 4140
rect 344986 4100 383660 4128
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 18598 4060 18604 4072
rect 14792 4032 18604 4060
rect 14792 4020 14798 4032
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 46658 4020 46664 4072
rect 46716 4060 46722 4072
rect 132865 4063 132923 4069
rect 132865 4060 132877 4063
rect 46716 4032 132877 4060
rect 46716 4020 46722 4032
rect 132865 4029 132877 4032
rect 132911 4029 132923 4063
rect 132865 4023 132923 4029
rect 132954 4020 132960 4072
rect 133012 4060 133018 4072
rect 133782 4060 133788 4072
rect 133012 4032 133788 4060
rect 133012 4020 133018 4032
rect 133782 4020 133788 4032
rect 133840 4020 133846 4072
rect 134150 4020 134156 4072
rect 134208 4060 134214 4072
rect 135162 4060 135168 4072
rect 134208 4032 135168 4060
rect 134208 4020 134214 4032
rect 135162 4020 135168 4032
rect 135220 4020 135226 4072
rect 280062 4020 280068 4072
rect 280120 4060 280126 4072
rect 344986 4060 345014 4100
rect 383654 4088 383660 4100
rect 383712 4088 383718 4140
rect 387150 4088 387156 4140
rect 387208 4128 387214 4140
rect 461210 4128 461216 4140
rect 387208 4100 461216 4128
rect 387208 4088 387214 4100
rect 461210 4088 461216 4100
rect 461268 4088 461274 4140
rect 461305 4131 461363 4137
rect 461305 4097 461317 4131
rect 461351 4128 461363 4131
rect 468018 4128 468024 4140
rect 461351 4100 468024 4128
rect 461351 4097 461363 4100
rect 461305 4091 461363 4097
rect 468018 4088 468024 4100
rect 468076 4088 468082 4140
rect 509329 4131 509387 4137
rect 509329 4128 509341 4131
rect 499546 4100 509341 4128
rect 280120 4032 345014 4060
rect 280120 4020 280126 4032
rect 383562 4020 383568 4072
rect 383620 4060 383626 4072
rect 461029 4063 461087 4069
rect 461029 4060 461041 4063
rect 383620 4032 461041 4060
rect 383620 4020 383626 4032
rect 461029 4029 461041 4032
rect 461075 4029 461087 4063
rect 461029 4023 461087 4029
rect 461118 4020 461124 4072
rect 461176 4060 461182 4072
rect 462406 4060 462412 4072
rect 461176 4032 462412 4060
rect 461176 4020 461182 4032
rect 462406 4020 462412 4032
rect 462464 4020 462470 4072
rect 462501 4063 462559 4069
rect 462501 4029 462513 4063
rect 462547 4060 462559 4063
rect 469214 4060 469220 4072
rect 462547 4032 469220 4060
rect 462547 4029 462559 4032
rect 462501 4023 462559 4029
rect 469214 4020 469220 4032
rect 469272 4020 469278 4072
rect 470686 4020 470692 4072
rect 470744 4060 470750 4072
rect 499546 4060 499574 4100
rect 509329 4097 509341 4100
rect 509375 4097 509387 4131
rect 509329 4091 509387 4097
rect 510522 4088 510528 4140
rect 510580 4128 510586 4140
rect 513929 4131 513987 4137
rect 513929 4128 513941 4131
rect 510580 4100 513941 4128
rect 510580 4088 510586 4100
rect 513929 4097 513941 4100
rect 513975 4097 513987 4131
rect 513929 4091 513987 4097
rect 514021 4131 514079 4137
rect 514021 4097 514033 4131
rect 514067 4128 514079 4131
rect 553762 4128 553768 4140
rect 514067 4100 553768 4128
rect 514067 4097 514079 4100
rect 514021 4091 514079 4097
rect 553762 4088 553768 4100
rect 553820 4088 553826 4140
rect 470744 4032 499574 4060
rect 470744 4020 470750 4032
rect 509142 4020 509148 4072
rect 509200 4060 509206 4072
rect 557350 4060 557356 4072
rect 509200 4032 557356 4060
rect 509200 4020 509206 4032
rect 557350 4020 557356 4032
rect 557408 4020 557414 4072
rect 43070 3952 43076 4004
rect 43128 3992 43134 4004
rect 138106 3992 138112 4004
rect 43128 3964 138112 3992
rect 43128 3952 43134 3964
rect 138106 3952 138112 3964
rect 138164 3952 138170 4004
rect 157794 3952 157800 4004
rect 157852 3992 157858 4004
rect 173894 3992 173900 4004
rect 157852 3964 173900 3992
rect 157852 3952 157858 3964
rect 173894 3952 173900 3964
rect 173952 3952 173958 4004
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 335998 3992 336004 4004
rect 333940 3964 336004 3992
rect 333940 3952 333946 3964
rect 335998 3952 336004 3964
rect 336056 3952 336062 4004
rect 379974 3952 379980 4004
rect 380032 3992 380038 4004
rect 460566 3992 460572 4004
rect 380032 3964 460572 3992
rect 380032 3952 380038 3964
rect 460566 3952 460572 3964
rect 460624 3952 460630 4004
rect 460842 3952 460848 4004
rect 460900 3992 460906 4004
rect 483198 3992 483204 4004
rect 460900 3964 483204 3992
rect 460900 3952 460906 3964
rect 483198 3952 483204 3964
rect 483256 3952 483262 4004
rect 489178 3952 489184 4004
rect 489236 3992 489242 4004
rect 492306 3992 492312 4004
rect 489236 3964 492312 3992
rect 489236 3952 489242 3964
rect 492306 3952 492312 3964
rect 492364 3952 492370 4004
rect 498010 3952 498016 4004
rect 498068 3992 498074 4004
rect 504453 3995 504511 4001
rect 504453 3992 504465 3995
rect 498068 3964 504465 3992
rect 498068 3952 498074 3964
rect 504453 3961 504465 3964
rect 504499 3961 504511 3995
rect 504453 3955 504511 3961
rect 509237 3995 509295 4001
rect 509237 3961 509249 3995
rect 509283 3992 509295 3995
rect 515950 3992 515956 4004
rect 509283 3964 515956 3992
rect 509283 3961 509295 3964
rect 509237 3955 509295 3961
rect 515950 3952 515956 3964
rect 516008 3952 516014 4004
rect 516137 3995 516195 4001
rect 516137 3961 516149 3995
rect 516183 3992 516195 3995
rect 560846 3992 560852 4004
rect 516183 3964 560852 3992
rect 516183 3961 516195 3964
rect 516137 3955 516195 3961
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 39574 3884 39580 3936
rect 39632 3924 39638 3936
rect 138014 3924 138020 3936
rect 39632 3896 138020 3924
rect 39632 3884 39638 3896
rect 138014 3884 138020 3896
rect 138072 3884 138078 3936
rect 154206 3884 154212 3936
rect 154264 3924 154270 3936
rect 172606 3924 172612 3936
rect 154264 3896 172612 3924
rect 154264 3884 154270 3896
rect 172606 3884 172612 3896
rect 172664 3884 172670 3936
rect 186038 3884 186044 3936
rect 186096 3924 186102 3936
rect 203886 3924 203892 3936
rect 186096 3896 203892 3924
rect 186096 3884 186102 3896
rect 203886 3884 203892 3896
rect 203944 3884 203950 3936
rect 276014 3884 276020 3936
rect 276072 3924 276078 3936
rect 277302 3924 277308 3936
rect 276072 3896 277308 3924
rect 276072 3884 276078 3896
rect 277302 3884 277308 3896
rect 277360 3884 277366 3936
rect 376478 3884 376484 3936
rect 376536 3924 376542 3936
rect 451277 3927 451335 3933
rect 451277 3924 451289 3927
rect 376536 3896 451289 3924
rect 376536 3884 376542 3896
rect 451277 3893 451289 3896
rect 451323 3893 451335 3927
rect 451277 3887 451335 3893
rect 451366 3884 451372 3936
rect 451424 3924 451430 3936
rect 455417 3927 455475 3933
rect 455417 3924 455429 3927
rect 451424 3896 455429 3924
rect 451424 3884 451430 3896
rect 455417 3893 455429 3896
rect 455463 3893 455475 3927
rect 455417 3887 455475 3893
rect 455506 3884 455512 3936
rect 455564 3924 455570 3936
rect 460658 3924 460664 3936
rect 455564 3896 460664 3924
rect 455564 3884 455570 3896
rect 460658 3884 460664 3896
rect 460716 3884 460722 3936
rect 460753 3927 460811 3933
rect 460753 3893 460765 3927
rect 460799 3924 460811 3927
rect 480622 3924 480628 3936
rect 460799 3896 480628 3924
rect 460799 3893 460811 3896
rect 460753 3887 460811 3893
rect 480622 3884 480628 3896
rect 480680 3884 480686 3936
rect 496722 3884 496728 3936
rect 496780 3924 496786 3936
rect 507670 3924 507676 3936
rect 496780 3896 507676 3924
rect 496780 3884 496786 3896
rect 507670 3884 507676 3896
rect 507728 3884 507734 3936
rect 509050 3884 509056 3936
rect 509108 3924 509114 3936
rect 514021 3927 514079 3933
rect 514021 3924 514033 3927
rect 509108 3896 514033 3924
rect 509108 3884 509114 3896
rect 514021 3893 514033 3896
rect 514067 3893 514079 3927
rect 514021 3887 514079 3893
rect 514113 3927 514171 3933
rect 514113 3893 514125 3927
rect 514159 3924 514171 3927
rect 564434 3924 564440 3936
rect 514159 3896 564440 3924
rect 514159 3893 514171 3896
rect 514113 3887 514171 3893
rect 564434 3884 564440 3896
rect 564492 3884 564498 3936
rect 1104 3760 582820 3856
rect 35986 3680 35992 3732
rect 36044 3720 36050 3732
rect 116305 3723 116363 3729
rect 116305 3720 116317 3723
rect 36044 3692 116317 3720
rect 36044 3680 36050 3692
rect 116305 3689 116317 3692
rect 116351 3689 116363 3723
rect 116305 3683 116363 3689
rect 116394 3680 116400 3732
rect 116452 3720 116458 3732
rect 117222 3720 117228 3732
rect 116452 3692 117228 3720
rect 116452 3680 116458 3692
rect 117222 3680 117228 3692
rect 117280 3680 117286 3732
rect 117590 3680 117596 3732
rect 117648 3720 117654 3732
rect 124585 3723 124643 3729
rect 124585 3720 124597 3723
rect 117648 3692 124597 3720
rect 117648 3680 117654 3692
rect 124585 3689 124597 3692
rect 124631 3689 124643 3723
rect 124585 3683 124643 3689
rect 124674 3680 124680 3732
rect 124732 3720 124738 3732
rect 158714 3720 158720 3732
rect 124732 3692 158720 3720
rect 124732 3680 124738 3692
rect 158714 3680 158720 3692
rect 158772 3680 158778 3732
rect 168374 3680 168380 3732
rect 168432 3720 168438 3732
rect 176010 3720 176016 3732
rect 168432 3692 176016 3720
rect 168432 3680 168438 3692
rect 176010 3680 176016 3692
rect 176068 3680 176074 3732
rect 187602 3680 187608 3732
rect 187660 3720 187666 3732
rect 207382 3720 207388 3732
rect 187660 3692 207388 3720
rect 187660 3680 187666 3692
rect 207382 3680 207388 3692
rect 207440 3680 207446 3732
rect 226334 3680 226340 3732
rect 226392 3720 226398 3732
rect 227530 3720 227536 3732
rect 226392 3692 227536 3720
rect 226392 3680 226398 3692
rect 227530 3680 227536 3692
rect 227588 3680 227594 3732
rect 251174 3680 251180 3732
rect 251232 3720 251238 3732
rect 252370 3720 252376 3732
rect 251232 3692 252376 3720
rect 251232 3680 251238 3692
rect 252370 3680 252376 3692
rect 252428 3680 252434 3732
rect 319714 3680 319720 3732
rect 319772 3720 319778 3732
rect 320818 3720 320824 3732
rect 319772 3692 320824 3720
rect 319772 3680 319778 3692
rect 320818 3680 320824 3692
rect 320876 3680 320882 3732
rect 358722 3680 358728 3732
rect 358780 3720 358786 3732
rect 451274 3720 451280 3732
rect 358780 3692 451280 3720
rect 358780 3680 358786 3692
rect 451274 3680 451280 3692
rect 451332 3680 451338 3732
rect 451369 3723 451427 3729
rect 451369 3689 451381 3723
rect 451415 3720 451427 3723
rect 454402 3720 454408 3732
rect 451415 3692 454408 3720
rect 451415 3689 451427 3692
rect 451369 3683 451427 3689
rect 454402 3680 454408 3692
rect 454460 3680 454466 3732
rect 454494 3680 454500 3732
rect 454552 3720 454558 3732
rect 455322 3720 455328 3732
rect 454552 3692 455328 3720
rect 454552 3680 454558 3692
rect 455322 3680 455328 3692
rect 455380 3680 455386 3732
rect 455417 3723 455475 3729
rect 455417 3689 455429 3723
rect 455463 3720 455475 3723
rect 477678 3720 477684 3732
rect 455463 3692 477684 3720
rect 455463 3689 455475 3692
rect 455417 3683 455475 3689
rect 477678 3680 477684 3692
rect 477736 3680 477742 3732
rect 495342 3680 495348 3732
rect 495400 3720 495406 3732
rect 500586 3720 500592 3732
rect 495400 3692 500592 3720
rect 495400 3680 495406 3692
rect 500586 3680 500592 3692
rect 500644 3680 500650 3732
rect 511258 3720 511264 3732
rect 504376 3692 511264 3720
rect 32490 3612 32496 3664
rect 32548 3652 32554 3664
rect 127621 3655 127679 3661
rect 127621 3652 127633 3655
rect 32548 3624 127633 3652
rect 32548 3612 32554 3624
rect 127621 3621 127633 3624
rect 127667 3621 127679 3655
rect 127621 3615 127679 3621
rect 127713 3655 127771 3661
rect 127713 3621 127725 3655
rect 127759 3652 127771 3655
rect 128541 3655 128599 3661
rect 127759 3624 128492 3652
rect 127759 3621 127771 3624
rect 127713 3615 127771 3621
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 14458 3584 14464 3596
rect 8812 3556 14464 3584
rect 8812 3544 8818 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 19978 3584 19984 3596
rect 15988 3556 19984 3584
rect 15988 3544 15994 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28902 3584 28908 3596
rect 27764 3556 28908 3584
rect 27764 3544 27770 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 31294 3544 31300 3596
rect 31352 3584 31358 3596
rect 32398 3584 32404 3596
rect 31352 3556 32404 3584
rect 31352 3544 31358 3556
rect 32398 3544 32404 3556
rect 32456 3544 32462 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34517 3587 34575 3593
rect 34517 3553 34529 3587
rect 34563 3584 34575 3587
rect 128464 3584 128492 3624
rect 128541 3621 128553 3655
rect 128587 3652 128599 3655
rect 136634 3652 136640 3664
rect 128587 3624 136640 3652
rect 128587 3621 128599 3624
rect 128541 3615 128599 3621
rect 136634 3612 136640 3624
rect 136692 3612 136698 3664
rect 158806 3652 158812 3664
rect 136744 3624 158812 3652
rect 133966 3584 133972 3596
rect 34563 3556 128400 3584
rect 128464 3556 133972 3584
rect 34563 3553 34575 3556
rect 34517 3547 34575 3553
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24268 3488 123432 3516
rect 24268 3476 24274 3488
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 10318 3448 10324 3460
rect 7708 3420 10324 3448
rect 7708 3408 7714 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 123297 3451 123355 3457
rect 123297 3448 123309 3451
rect 19484 3420 123309 3448
rect 19484 3408 19490 3420
rect 123297 3417 123309 3420
rect 123343 3417 123355 3451
rect 123404 3448 123432 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124585 3519 124643 3525
rect 124585 3485 124597 3519
rect 124631 3516 124643 3519
rect 126885 3519 126943 3525
rect 126885 3516 126897 3519
rect 124631 3488 126897 3516
rect 124631 3485 124643 3488
rect 124585 3479 124643 3485
rect 126885 3485 126897 3488
rect 126931 3485 126943 3519
rect 126885 3479 126943 3485
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128262 3516 128268 3528
rect 127032 3488 128268 3516
rect 127032 3476 127038 3488
rect 128262 3476 128268 3488
rect 128320 3476 128326 3528
rect 128372 3516 128400 3556
rect 133966 3544 133972 3556
rect 134024 3544 134030 3596
rect 134058 3544 134064 3596
rect 134116 3584 134122 3596
rect 136744 3584 136772 3624
rect 158806 3612 158812 3624
rect 158864 3612 158870 3664
rect 160094 3612 160100 3664
rect 160152 3652 160158 3664
rect 405734 3652 405740 3664
rect 160152 3624 405740 3652
rect 160152 3612 160158 3624
rect 405734 3612 405740 3624
rect 405792 3612 405798 3664
rect 415486 3612 415492 3664
rect 415544 3652 415550 3664
rect 416682 3652 416688 3664
rect 415544 3624 416688 3652
rect 415544 3612 415550 3624
rect 416682 3612 416688 3624
rect 416740 3612 416746 3664
rect 422570 3612 422576 3664
rect 422628 3652 422634 3664
rect 423582 3652 423588 3664
rect 422628 3624 423588 3652
rect 422628 3612 422634 3624
rect 423582 3612 423588 3624
rect 423640 3612 423646 3664
rect 426069 3655 426127 3661
rect 426069 3621 426081 3655
rect 426115 3652 426127 3655
rect 473538 3652 473544 3664
rect 426115 3624 473544 3652
rect 426115 3621 426127 3624
rect 426069 3615 426127 3621
rect 473538 3612 473544 3624
rect 473596 3612 473602 3664
rect 498102 3612 498108 3664
rect 498160 3652 498166 3664
rect 504376 3652 504404 3692
rect 511258 3680 511264 3692
rect 511316 3680 511322 3732
rect 511810 3680 511816 3732
rect 511868 3720 511874 3732
rect 514113 3723 514171 3729
rect 514113 3720 514125 3723
rect 511868 3692 514125 3720
rect 511868 3680 511874 3692
rect 514113 3689 514125 3692
rect 514159 3689 514171 3723
rect 514113 3683 514171 3689
rect 514205 3723 514263 3729
rect 514205 3689 514217 3723
rect 514251 3720 514263 3723
rect 516137 3723 516195 3729
rect 516137 3720 516149 3723
rect 514251 3692 516149 3720
rect 514251 3689 514263 3692
rect 514205 3683 514263 3689
rect 516137 3689 516149 3692
rect 516183 3689 516195 3723
rect 516137 3683 516195 3689
rect 516226 3680 516232 3732
rect 516284 3720 516290 3732
rect 516284 3692 518572 3720
rect 516284 3680 516290 3692
rect 498160 3624 504404 3652
rect 504453 3655 504511 3661
rect 498160 3612 498166 3624
rect 504453 3621 504465 3655
rect 504499 3652 504511 3655
rect 514754 3652 514760 3664
rect 504499 3624 514760 3652
rect 504499 3621 504511 3624
rect 504453 3615 504511 3621
rect 514754 3612 514760 3624
rect 514812 3612 514818 3664
rect 516042 3612 516048 3664
rect 516100 3652 516106 3664
rect 518544 3652 518572 3692
rect 518618 3680 518624 3732
rect 518676 3720 518682 3732
rect 568022 3720 568028 3732
rect 518676 3692 568028 3720
rect 518676 3680 518682 3692
rect 568022 3680 568028 3692
rect 568080 3680 568086 3732
rect 571518 3652 571524 3664
rect 516100 3624 518480 3652
rect 518544 3624 571524 3652
rect 516100 3612 516106 3624
rect 139394 3584 139400 3596
rect 134116 3556 136772 3584
rect 137986 3556 139400 3584
rect 134116 3544 134122 3556
rect 128449 3519 128507 3525
rect 128449 3516 128461 3519
rect 128372 3488 128461 3516
rect 128449 3485 128461 3488
rect 128495 3485 128507 3519
rect 132773 3519 132831 3525
rect 132773 3516 132785 3519
rect 128449 3479 128507 3485
rect 128556 3488 132785 3516
rect 127529 3451 127587 3457
rect 127529 3448 127541 3451
rect 123404 3420 127541 3448
rect 123297 3411 123355 3417
rect 127529 3417 127541 3420
rect 127575 3417 127587 3451
rect 127529 3411 127587 3417
rect 127621 3451 127679 3457
rect 127621 3417 127633 3451
rect 127667 3448 127679 3451
rect 128556 3448 128584 3488
rect 132773 3485 132785 3488
rect 132819 3485 132831 3519
rect 132773 3479 132831 3485
rect 132865 3519 132923 3525
rect 132865 3485 132877 3519
rect 132911 3516 132923 3519
rect 137986 3516 138014 3556
rect 139394 3544 139400 3556
rect 139452 3544 139458 3596
rect 143534 3544 143540 3596
rect 143592 3584 143598 3596
rect 144730 3584 144736 3596
rect 143592 3556 144736 3584
rect 143592 3544 143598 3556
rect 144730 3544 144736 3556
rect 144788 3544 144794 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 405826 3584 405832 3596
rect 156656 3556 405832 3584
rect 156656 3544 156662 3556
rect 405826 3544 405832 3556
rect 405884 3544 405890 3596
rect 411898 3544 411904 3596
rect 411956 3584 411962 3596
rect 470778 3584 470784 3596
rect 411956 3556 470784 3584
rect 411956 3544 411962 3556
rect 470778 3544 470784 3556
rect 470836 3544 470842 3596
rect 485038 3544 485044 3596
rect 485096 3544 485102 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 491202 3584 491208 3596
rect 489972 3556 491208 3584
rect 489972 3544 489978 3556
rect 491202 3544 491208 3556
rect 491260 3544 491266 3596
rect 499298 3544 499304 3596
rect 499356 3584 499362 3596
rect 518342 3584 518348 3596
rect 499356 3556 518348 3584
rect 499356 3544 499362 3556
rect 518342 3544 518348 3556
rect 518400 3544 518406 3596
rect 518452 3584 518480 3624
rect 571518 3612 571524 3624
rect 571576 3612 571582 3664
rect 523589 3587 523647 3593
rect 523589 3584 523601 3587
rect 518452 3556 523601 3584
rect 523589 3553 523601 3556
rect 523635 3553 523647 3587
rect 575106 3584 575112 3596
rect 523589 3547 523647 3553
rect 523696 3556 575112 3584
rect 132911 3488 138014 3516
rect 132911 3485 132923 3488
rect 132865 3479 132923 3485
rect 138842 3476 138848 3528
rect 138900 3516 138906 3528
rect 139302 3516 139308 3528
rect 138900 3488 139308 3516
rect 138900 3476 138906 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151722 3516 151728 3528
rect 150676 3488 151728 3516
rect 150676 3476 150682 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 155402 3476 155408 3528
rect 155460 3516 155466 3528
rect 155862 3516 155868 3528
rect 155460 3488 155868 3516
rect 155460 3476 155466 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156969 3519 157027 3525
rect 156969 3485 156981 3519
rect 157015 3516 157027 3519
rect 404354 3516 404360 3528
rect 157015 3488 404360 3516
rect 157015 3485 157027 3488
rect 156969 3479 157027 3485
rect 404354 3476 404360 3488
rect 404412 3476 404418 3528
rect 408402 3476 408408 3528
rect 408460 3516 408466 3528
rect 470594 3516 470600 3528
rect 408460 3488 470600 3516
rect 408460 3476 408466 3488
rect 470594 3476 470600 3488
rect 470652 3476 470658 3528
rect 479334 3476 479340 3528
rect 479392 3516 479398 3528
rect 480162 3516 480168 3528
rect 479392 3488 480168 3516
rect 479392 3476 479398 3488
rect 480162 3476 480168 3488
rect 480220 3476 480226 3528
rect 127667 3420 128584 3448
rect 128633 3451 128691 3457
rect 127667 3417 127679 3420
rect 127621 3411 127679 3417
rect 128633 3417 128645 3451
rect 128679 3448 128691 3451
rect 135254 3448 135260 3460
rect 128679 3420 135260 3448
rect 128679 3417 128691 3420
rect 128633 3411 128691 3417
rect 135254 3408 135260 3420
rect 135312 3408 135318 3460
rect 149514 3408 149520 3460
rect 149572 3448 149578 3460
rect 158533 3451 158591 3457
rect 158533 3448 158545 3451
rect 149572 3420 158545 3448
rect 149572 3408 149578 3420
rect 158533 3417 158545 3420
rect 158579 3417 158591 3451
rect 158533 3411 158591 3417
rect 158717 3451 158775 3457
rect 158717 3417 158729 3451
rect 158763 3448 158775 3451
rect 402974 3448 402980 3460
rect 158763 3420 402980 3448
rect 158763 3417 158775 3420
rect 158717 3411 158775 3417
rect 402974 3408 402980 3420
rect 403032 3408 403038 3460
rect 404814 3408 404820 3460
rect 404872 3448 404878 3460
rect 461489 3451 461547 3457
rect 461489 3448 461501 3451
rect 404872 3420 461501 3448
rect 404872 3408 404878 3420
rect 461489 3417 461501 3420
rect 461535 3417 461547 3451
rect 461489 3411 461547 3417
rect 461578 3408 461584 3460
rect 461636 3448 461642 3460
rect 462222 3448 462228 3460
rect 461636 3420 462228 3448
rect 461636 3408 461642 3420
rect 462222 3408 462228 3420
rect 462280 3408 462286 3460
rect 462314 3408 462320 3460
rect 462372 3448 462378 3460
rect 467926 3448 467932 3460
rect 462372 3420 467932 3448
rect 462372 3408 462378 3420
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 468662 3408 468668 3460
rect 468720 3448 468726 3460
rect 469122 3448 469128 3460
rect 468720 3420 469128 3448
rect 468720 3408 468726 3420
rect 469122 3408 469128 3420
rect 469180 3408 469186 3460
rect 485056 3448 485084 3544
rect 486418 3476 486424 3528
rect 486476 3516 486482 3528
rect 487062 3516 487068 3528
rect 486476 3488 487068 3516
rect 486476 3476 486482 3488
rect 487062 3476 487068 3488
rect 487120 3476 487126 3528
rect 487798 3476 487804 3528
rect 487856 3516 487862 3528
rect 487856 3488 493824 3516
rect 487856 3476 487862 3488
rect 493796 3448 493824 3488
rect 493962 3476 493968 3528
rect 494020 3516 494026 3528
rect 497090 3516 497096 3528
rect 494020 3488 497096 3516
rect 494020 3476 494026 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 500770 3476 500776 3528
rect 500828 3516 500834 3528
rect 521838 3516 521844 3528
rect 500828 3488 521844 3516
rect 500828 3476 500834 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 521933 3519 521991 3525
rect 521933 3485 521945 3519
rect 521979 3516 521991 3519
rect 523696 3516 523724 3556
rect 575106 3544 575112 3556
rect 575164 3544 575170 3596
rect 521979 3488 523724 3516
rect 523773 3519 523831 3525
rect 521979 3485 521991 3488
rect 521933 3479 521991 3485
rect 523773 3485 523785 3519
rect 523819 3516 523831 3519
rect 579798 3516 579804 3528
rect 523819 3488 579804 3516
rect 523819 3485 523831 3488
rect 523773 3479 523831 3485
rect 579798 3476 579804 3488
rect 579856 3476 579862 3528
rect 495894 3448 495900 3460
rect 485056 3420 489914 3448
rect 493796 3420 495900 3448
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 34517 3383 34575 3389
rect 34517 3380 34529 3383
rect 28960 3352 34529 3380
rect 28960 3340 28966 3352
rect 34517 3349 34529 3352
rect 34563 3349 34575 3383
rect 34517 3343 34575 3349
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42702 3380 42708 3392
rect 41932 3352 42708 3380
rect 41932 3340 41938 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45370 3380 45376 3392
rect 44324 3352 45376 3380
rect 44324 3340 44330 3352
rect 45370 3340 45376 3352
rect 45428 3340 45434 3392
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 53650 3380 53656 3392
rect 52604 3352 53656 3380
rect 52604 3340 52610 3352
rect 53650 3340 53656 3352
rect 53708 3340 53714 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 57882 3380 57888 3392
rect 57296 3352 57888 3380
rect 57296 3340 57302 3352
rect 57882 3340 57888 3352
rect 57940 3340 57946 3392
rect 58434 3340 58440 3392
rect 58492 3380 58498 3392
rect 59262 3380 59268 3392
rect 58492 3352 59268 3380
rect 58492 3340 58498 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 60642 3380 60648 3392
rect 59688 3352 60648 3380
rect 59688 3340 59694 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 60826 3340 60832 3392
rect 60884 3380 60890 3392
rect 61930 3380 61936 3392
rect 60884 3352 61936 3380
rect 60884 3340 60890 3352
rect 61930 3340 61936 3352
rect 61988 3340 61994 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 68922 3380 68928 3392
rect 67968 3352 68928 3380
rect 67968 3340 67974 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 75822 3380 75828 3392
rect 75052 3352 75828 3380
rect 75052 3340 75058 3352
rect 75822 3340 75828 3352
rect 75880 3340 75886 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 82078 3340 82084 3392
rect 82136 3380 82142 3392
rect 82722 3380 82728 3392
rect 82136 3352 82728 3380
rect 82136 3340 82142 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 85482 3380 85488 3392
rect 84528 3352 85488 3380
rect 84528 3340 84534 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 92382 3380 92388 3392
rect 91612 3352 92388 3380
rect 91612 3340 91618 3352
rect 92382 3340 92388 3352
rect 92440 3340 92446 3392
rect 92477 3383 92535 3389
rect 92477 3349 92489 3383
rect 92523 3380 92535 3383
rect 150526 3380 150532 3392
rect 92523 3352 150532 3380
rect 92523 3349 92535 3352
rect 92477 3343 92535 3349
rect 150526 3340 150532 3352
rect 150584 3340 150590 3392
rect 153010 3340 153016 3392
rect 153068 3380 153074 3392
rect 156969 3383 157027 3389
rect 156969 3380 156981 3383
rect 153068 3352 156981 3380
rect 153068 3340 153074 3352
rect 156969 3349 156981 3352
rect 157015 3349 157027 3383
rect 156969 3343 157027 3349
rect 167178 3340 167184 3392
rect 167236 3380 167242 3392
rect 168282 3380 168288 3392
rect 167236 3352 168288 3380
rect 167236 3340 167242 3352
rect 168282 3340 168288 3352
rect 168340 3340 168346 3392
rect 174262 3340 174268 3392
rect 174320 3380 174326 3392
rect 175182 3380 175188 3392
rect 174320 3352 175188 3380
rect 174320 3340 174326 3352
rect 175182 3340 175188 3352
rect 175240 3340 175246 3392
rect 175458 3340 175464 3392
rect 175516 3380 175522 3392
rect 178126 3380 178132 3392
rect 175516 3352 178132 3380
rect 175516 3340 175522 3352
rect 178126 3340 178132 3352
rect 178184 3340 178190 3392
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 181990 3380 181996 3392
rect 181496 3352 181996 3380
rect 181496 3340 181502 3352
rect 181990 3340 181996 3352
rect 182048 3340 182054 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186130 3380 186136 3392
rect 184992 3352 186136 3380
rect 184992 3340 184998 3352
rect 186130 3340 186136 3352
rect 186188 3340 186194 3392
rect 206186 3340 206192 3392
rect 206244 3380 206250 3392
rect 206922 3380 206928 3392
rect 206244 3352 206928 3380
rect 206244 3340 206250 3352
rect 206922 3340 206928 3352
rect 206980 3340 206986 3392
rect 209774 3340 209780 3392
rect 209832 3380 209838 3392
rect 211062 3380 211068 3392
rect 209832 3352 211068 3380
rect 209832 3340 209838 3352
rect 211062 3340 211068 3352
rect 211120 3340 211126 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 216858 3340 216864 3392
rect 216916 3380 216922 3392
rect 217962 3380 217968 3392
rect 216916 3352 217968 3380
rect 216916 3340 216922 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 222746 3340 222752 3392
rect 222804 3380 222810 3392
rect 223298 3380 223304 3392
rect 222804 3352 223304 3380
rect 222804 3340 222810 3352
rect 223298 3340 223304 3352
rect 223356 3340 223362 3392
rect 223942 3340 223948 3392
rect 224000 3380 224006 3392
rect 224770 3380 224776 3392
rect 224000 3352 224776 3380
rect 224000 3340 224006 3352
rect 224770 3340 224776 3352
rect 224828 3340 224834 3392
rect 229830 3340 229836 3392
rect 229888 3380 229894 3392
rect 230382 3380 230388 3392
rect 229888 3352 230388 3380
rect 229888 3340 229894 3352
rect 230382 3340 230388 3352
rect 230440 3340 230446 3392
rect 231026 3340 231032 3392
rect 231084 3380 231090 3392
rect 231670 3380 231676 3392
rect 231084 3352 231676 3380
rect 231084 3340 231090 3352
rect 231670 3340 231676 3352
rect 231728 3340 231734 3392
rect 233418 3340 233424 3392
rect 233476 3380 233482 3392
rect 234430 3380 234436 3392
rect 233476 3352 234436 3380
rect 233476 3340 233482 3352
rect 234430 3340 234436 3352
rect 234488 3340 234494 3392
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235810 3380 235816 3392
rect 234672 3352 235816 3380
rect 234672 3340 234678 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 238110 3340 238116 3392
rect 238168 3380 238174 3392
rect 238662 3380 238668 3392
rect 238168 3352 238668 3380
rect 238168 3340 238174 3352
rect 238662 3340 238668 3352
rect 238720 3340 238726 3392
rect 240502 3340 240508 3392
rect 240560 3380 240566 3392
rect 241422 3380 241428 3392
rect 240560 3352 241428 3380
rect 240560 3340 240566 3352
rect 241422 3340 241428 3352
rect 241480 3340 241486 3392
rect 241698 3340 241704 3392
rect 241756 3380 241762 3392
rect 242618 3380 242624 3392
rect 241756 3352 242624 3380
rect 241756 3340 241762 3352
rect 242618 3340 242624 3352
rect 242676 3340 242682 3392
rect 247586 3340 247592 3392
rect 247644 3380 247650 3392
rect 248138 3380 248144 3392
rect 247644 3352 248144 3380
rect 247644 3340 247650 3352
rect 248138 3340 248144 3352
rect 248196 3340 248202 3392
rect 248782 3340 248788 3392
rect 248840 3380 248846 3392
rect 249610 3380 249616 3392
rect 248840 3352 249616 3380
rect 248840 3340 248846 3352
rect 249610 3340 249616 3352
rect 249668 3340 249674 3392
rect 254670 3340 254676 3392
rect 254728 3380 254734 3392
rect 255222 3380 255228 3392
rect 254728 3352 255228 3380
rect 254728 3340 254734 3352
rect 255222 3340 255228 3352
rect 255280 3340 255286 3392
rect 255866 3340 255872 3392
rect 255924 3380 255930 3392
rect 256418 3380 256424 3392
rect 255924 3352 256424 3380
rect 255924 3340 255930 3352
rect 256418 3340 256424 3352
rect 256476 3340 256482 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260558 3380 260564 3392
rect 259512 3352 260564 3380
rect 259512 3340 259518 3352
rect 260558 3340 260564 3352
rect 260616 3340 260622 3392
rect 265342 3340 265348 3392
rect 265400 3380 265406 3392
rect 266078 3380 266084 3392
rect 265400 3352 266084 3380
rect 265400 3340 265406 3352
rect 266078 3340 266084 3352
rect 266136 3340 266142 3392
rect 266538 3340 266544 3392
rect 266596 3380 266602 3392
rect 267550 3380 267556 3392
rect 266596 3352 267556 3380
rect 266596 3340 266602 3352
rect 267550 3340 267556 3352
rect 267608 3340 267614 3392
rect 272426 3340 272432 3392
rect 272484 3380 272490 3392
rect 273070 3380 273076 3392
rect 272484 3352 273076 3380
rect 272484 3340 272490 3352
rect 273070 3340 273076 3352
rect 273128 3340 273134 3392
rect 312630 3340 312636 3392
rect 312688 3380 312694 3392
rect 313182 3380 313188 3392
rect 312688 3352 313188 3380
rect 312688 3340 312694 3352
rect 313182 3340 313188 3352
rect 313240 3340 313246 3392
rect 316218 3340 316224 3392
rect 316276 3380 316282 3392
rect 318058 3380 318064 3392
rect 316276 3352 318064 3380
rect 316276 3340 316282 3352
rect 318058 3340 318064 3352
rect 318116 3340 318122 3392
rect 323302 3340 323308 3392
rect 323360 3380 323366 3392
rect 324222 3380 324228 3392
rect 323360 3352 324228 3380
rect 323360 3340 323366 3352
rect 324222 3340 324228 3352
rect 324280 3340 324286 3392
rect 330386 3340 330392 3392
rect 330444 3380 330450 3392
rect 331122 3380 331128 3392
rect 330444 3352 331128 3380
rect 330444 3340 330450 3352
rect 331122 3340 331128 3352
rect 331180 3340 331186 3392
rect 335354 3340 335360 3392
rect 335412 3380 335418 3392
rect 336274 3380 336280 3392
rect 335412 3352 336280 3380
rect 335412 3340 335418 3352
rect 336274 3340 336280 3352
rect 336332 3340 336338 3392
rect 337470 3340 337476 3392
rect 337528 3380 337534 3392
rect 338758 3380 338764 3392
rect 337528 3352 338764 3380
rect 337528 3340 337534 3352
rect 338758 3340 338764 3352
rect 338816 3340 338822 3392
rect 348050 3340 348056 3392
rect 348108 3380 348114 3392
rect 349798 3380 349804 3392
rect 348108 3352 349804 3380
rect 348108 3340 348114 3352
rect 349798 3340 349804 3352
rect 349856 3340 349862 3392
rect 351638 3340 351644 3392
rect 351696 3380 351702 3392
rect 352558 3380 352564 3392
rect 351696 3352 352564 3380
rect 351696 3340 351702 3352
rect 352558 3340 352564 3352
rect 352616 3340 352622 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 460937 3383 460995 3389
rect 460937 3380 460949 3383
rect 390704 3352 460949 3380
rect 390704 3340 390710 3352
rect 460937 3349 460949 3352
rect 460983 3349 460995 3383
rect 460937 3343 460995 3349
rect 461029 3383 461087 3389
rect 461029 3349 461041 3383
rect 461075 3380 461087 3383
rect 463694 3380 463700 3392
rect 461075 3352 463700 3380
rect 461075 3349 461087 3352
rect 461029 3343 461087 3349
rect 463694 3340 463700 3352
rect 463752 3340 463758 3392
rect 489886 3380 489914 3420
rect 495894 3408 495900 3420
rect 495952 3408 495958 3460
rect 500862 3408 500868 3460
rect 500920 3448 500926 3460
rect 518897 3451 518955 3457
rect 518897 3448 518909 3451
rect 500920 3420 518909 3448
rect 500920 3408 500926 3420
rect 518897 3417 518909 3420
rect 518943 3417 518955 3451
rect 518897 3411 518955 3417
rect 518986 3408 518992 3460
rect 519044 3448 519050 3460
rect 583386 3448 583392 3460
rect 519044 3420 583392 3448
rect 519044 3408 519050 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 499390 3380 499396 3392
rect 489886 3352 499396 3380
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 507762 3340 507768 3392
rect 507820 3380 507826 3392
rect 550266 3380 550272 3392
rect 507820 3352 550272 3380
rect 507820 3340 507826 3352
rect 550266 3340 550272 3352
rect 550324 3340 550330 3392
rect 1104 3216 582820 3312
rect 89162 3136 89168 3188
rect 89220 3176 89226 3188
rect 92477 3179 92535 3185
rect 92477 3176 92489 3179
rect 89220 3148 92489 3176
rect 89220 3136 89226 3148
rect 92477 3145 92489 3148
rect 92523 3145 92535 3179
rect 92477 3139 92535 3145
rect 92750 3136 92756 3188
rect 92808 3176 92814 3188
rect 150434 3176 150440 3188
rect 92808 3148 150440 3176
rect 92808 3136 92814 3148
rect 150434 3136 150440 3148
rect 150492 3136 150498 3188
rect 171962 3136 171968 3188
rect 172020 3176 172026 3188
rect 175918 3176 175924 3188
rect 172020 3148 175924 3176
rect 172020 3136 172026 3148
rect 175918 3136 175924 3148
rect 175976 3136 175982 3188
rect 182082 3136 182088 3188
rect 182140 3176 182146 3188
rect 186130 3176 186136 3188
rect 182140 3148 186136 3176
rect 182140 3136 182146 3148
rect 186130 3136 186136 3148
rect 186188 3136 186194 3188
rect 199102 3136 199108 3188
rect 199160 3176 199166 3188
rect 199838 3176 199844 3188
rect 199160 3148 199844 3176
rect 199160 3136 199166 3148
rect 199838 3136 199844 3148
rect 199896 3136 199902 3188
rect 322106 3136 322112 3188
rect 322164 3176 322170 3188
rect 322842 3176 322848 3188
rect 322164 3148 322848 3176
rect 322164 3136 322170 3148
rect 322842 3136 322848 3148
rect 322900 3136 322906 3188
rect 390554 3136 390560 3188
rect 390612 3176 390618 3188
rect 391842 3176 391848 3188
rect 390612 3148 391848 3176
rect 390612 3136 390618 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 394234 3136 394240 3188
rect 394292 3176 394298 3188
rect 394292 3148 461164 3176
rect 394292 3136 394298 3148
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 17862 3108 17868 3120
rect 17092 3080 17868 3108
rect 17092 3068 17098 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 99834 3068 99840 3120
rect 99892 3108 99898 3120
rect 153194 3108 153200 3120
rect 99892 3080 153200 3108
rect 99892 3068 99898 3080
rect 153194 3068 153200 3080
rect 153252 3068 153258 3120
rect 397730 3068 397736 3120
rect 397788 3108 397794 3120
rect 460842 3108 460848 3120
rect 397788 3080 460848 3108
rect 397788 3068 397794 3080
rect 460842 3068 460848 3080
rect 460900 3068 460906 3120
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 15838 3040 15844 3052
rect 13596 3012 15844 3040
rect 13596 3000 13602 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 103330 3000 103336 3052
rect 103388 3040 103394 3052
rect 153286 3040 153292 3052
rect 103388 3012 153292 3040
rect 103388 3000 103394 3012
rect 153286 3000 153292 3012
rect 153344 3000 153350 3052
rect 340966 3000 340972 3052
rect 341024 3040 341030 3052
rect 344278 3040 344284 3052
rect 341024 3012 344284 3040
rect 341024 3000 341030 3012
rect 344278 3000 344284 3012
rect 344336 3000 344342 3052
rect 355226 3000 355232 3052
rect 355284 3040 355290 3052
rect 358078 3040 358084 3052
rect 355284 3012 358084 3040
rect 355284 3000 355290 3012
rect 358078 3000 358084 3012
rect 358136 3000 358142 3052
rect 401318 3000 401324 3052
rect 401376 3040 401382 3052
rect 461029 3043 461087 3049
rect 461029 3040 461041 3043
rect 401376 3012 461041 3040
rect 401376 3000 401382 3012
rect 461029 3009 461041 3012
rect 461075 3009 461087 3043
rect 461136 3040 461164 3148
rect 461302 3136 461308 3188
rect 461360 3176 461366 3188
rect 465074 3176 465080 3188
rect 461360 3148 465080 3176
rect 461360 3136 461366 3148
rect 465074 3136 465080 3148
rect 465132 3136 465138 3188
rect 465166 3136 465172 3188
rect 465224 3176 465230 3188
rect 466362 3176 466368 3188
rect 465224 3148 466368 3176
rect 465224 3136 465230 3148
rect 466362 3136 466368 3148
rect 466420 3136 466426 3188
rect 472250 3136 472256 3188
rect 472308 3176 472314 3188
rect 473262 3176 473268 3188
rect 472308 3148 473268 3176
rect 472308 3136 472314 3148
rect 473262 3136 473268 3148
rect 473320 3136 473326 3188
rect 506382 3136 506388 3188
rect 506440 3176 506446 3188
rect 546678 3176 546684 3188
rect 506440 3148 546684 3176
rect 506440 3136 506446 3148
rect 546678 3136 546684 3148
rect 546736 3136 546742 3188
rect 461213 3111 461271 3117
rect 461213 3077 461225 3111
rect 461259 3108 461271 3111
rect 465350 3108 465356 3120
rect 461259 3080 465356 3108
rect 461259 3077 461271 3080
rect 461213 3071 461271 3077
rect 465350 3068 465356 3080
rect 465408 3068 465414 3120
rect 506290 3068 506296 3120
rect 506348 3108 506354 3120
rect 543182 3108 543188 3120
rect 506348 3080 543188 3108
rect 506348 3068 506354 3080
rect 543182 3068 543188 3080
rect 543240 3068 543246 3120
rect 466454 3040 466460 3052
rect 461136 3012 466460 3040
rect 461029 3003 461087 3009
rect 466454 3000 466460 3012
rect 466512 3000 466518 3052
rect 505002 3000 505008 3052
rect 505060 3040 505066 3052
rect 539594 3040 539600 3052
rect 505060 3012 539600 3040
rect 505060 3000 505066 3012
rect 539594 3000 539600 3012
rect 539652 3000 539658 3052
rect 105722 2932 105728 2984
rect 105780 2972 105786 2984
rect 106182 2972 106188 2984
rect 105780 2944 106188 2972
rect 105780 2932 105786 2944
rect 106182 2932 106188 2944
rect 106240 2932 106246 2984
rect 106918 2932 106924 2984
rect 106976 2972 106982 2984
rect 107562 2972 107568 2984
rect 106976 2944 107568 2972
rect 106976 2932 106982 2944
rect 107562 2932 107568 2944
rect 107620 2932 107626 2984
rect 109310 2932 109316 2984
rect 109368 2972 109374 2984
rect 110322 2972 110328 2984
rect 109368 2944 110328 2972
rect 109368 2932 109374 2944
rect 110322 2932 110328 2944
rect 110380 2932 110386 2984
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 155954 2972 155960 2984
rect 110564 2944 155960 2972
rect 110564 2932 110570 2944
rect 155954 2932 155960 2944
rect 156012 2932 156018 2984
rect 192018 2932 192024 2984
rect 192076 2972 192082 2984
rect 193030 2972 193036 2984
rect 192076 2944 193036 2972
rect 192076 2932 192082 2944
rect 193030 2932 193036 2944
rect 193088 2932 193094 2984
rect 258258 2932 258264 2984
rect 258316 2972 258322 2984
rect 259362 2972 259368 2984
rect 258316 2944 259368 2972
rect 258316 2932 258322 2944
rect 259362 2932 259368 2944
rect 259420 2932 259426 2984
rect 415486 2932 415492 2984
rect 415544 2972 415550 2984
rect 416590 2972 416596 2984
rect 415544 2944 416596 2972
rect 415544 2932 415550 2944
rect 416590 2932 416596 2944
rect 416648 2932 416654 2984
rect 418982 2932 418988 2984
rect 419040 2972 419046 2984
rect 426069 2975 426127 2981
rect 426069 2972 426081 2975
rect 419040 2944 426081 2972
rect 419040 2932 419046 2944
rect 426069 2941 426081 2944
rect 426115 2941 426127 2975
rect 426069 2935 426127 2941
rect 426158 2932 426164 2984
rect 426216 2972 426222 2984
rect 474826 2972 474832 2984
rect 426216 2944 474832 2972
rect 426216 2932 426222 2944
rect 474826 2932 474832 2944
rect 474884 2932 474890 2984
rect 503622 2932 503628 2984
rect 503680 2972 503686 2984
rect 536098 2972 536104 2984
rect 503680 2944 536104 2972
rect 503680 2932 503686 2944
rect 536098 2932 536104 2944
rect 536156 2932 536162 2984
rect 73798 2864 73804 2916
rect 73856 2904 73862 2916
rect 74442 2904 74448 2916
rect 73856 2876 74448 2904
rect 73856 2864 73862 2876
rect 74442 2864 74448 2876
rect 74500 2864 74506 2916
rect 114002 2864 114008 2916
rect 114060 2904 114066 2916
rect 156046 2904 156052 2916
rect 114060 2876 156052 2904
rect 114060 2864 114066 2876
rect 156046 2864 156052 2876
rect 156104 2864 156110 2916
rect 280706 2864 280712 2916
rect 280764 2904 280770 2916
rect 281442 2904 281448 2916
rect 280764 2876 281448 2904
rect 280764 2864 280770 2876
rect 281442 2864 281448 2876
rect 281500 2864 281506 2916
rect 429654 2864 429660 2916
rect 429712 2904 429718 2916
rect 476114 2904 476120 2916
rect 429712 2876 476120 2904
rect 429712 2864 429718 2876
rect 476114 2864 476120 2876
rect 476172 2864 476178 2916
rect 503530 2864 503536 2916
rect 503588 2904 503594 2916
rect 532510 2904 532516 2916
rect 503588 2876 532516 2904
rect 503588 2864 503594 2876
rect 532510 2864 532516 2876
rect 532568 2864 532574 2916
rect 116305 2839 116363 2845
rect 116305 2805 116317 2839
rect 116351 2836 116363 2839
rect 123205 2839 123263 2845
rect 123205 2836 123217 2839
rect 116351 2808 123217 2836
rect 116351 2805 116363 2808
rect 116305 2799 116363 2805
rect 123205 2805 123217 2808
rect 123251 2805 123263 2839
rect 123205 2799 123263 2805
rect 123297 2839 123355 2845
rect 123297 2805 123309 2839
rect 123343 2836 123355 2839
rect 128354 2836 128360 2848
rect 123343 2808 128360 2836
rect 123343 2805 123355 2808
rect 123297 2799 123355 2805
rect 128354 2796 128360 2808
rect 128412 2796 128418 2848
rect 128449 2839 128507 2845
rect 128449 2805 128461 2839
rect 128495 2836 128507 2839
rect 132218 2836 132224 2848
rect 128495 2808 132224 2836
rect 128495 2805 128507 2808
rect 128449 2799 128507 2805
rect 132218 2796 132224 2808
rect 132276 2796 132282 2848
rect 132313 2839 132371 2845
rect 132313 2805 132325 2839
rect 132359 2836 132371 2839
rect 157334 2836 157340 2848
rect 132359 2808 157340 2836
rect 132359 2805 132371 2808
rect 132313 2799 132371 2805
rect 157334 2796 157340 2808
rect 157392 2796 157398 2848
rect 433242 2796 433248 2848
rect 433300 2836 433306 2848
rect 436649 2839 436707 2845
rect 436649 2836 436661 2839
rect 433300 2808 436661 2836
rect 433300 2796 433306 2808
rect 436649 2805 436661 2808
rect 436695 2805 436707 2839
rect 436649 2799 436707 2805
rect 436738 2796 436744 2848
rect 436796 2836 436802 2848
rect 437382 2836 437388 2848
rect 436796 2808 437388 2836
rect 436796 2796 436802 2808
rect 437382 2796 437388 2808
rect 437440 2796 437446 2848
rect 437477 2839 437535 2845
rect 437477 2805 437489 2839
rect 437523 2836 437535 2839
rect 476206 2836 476212 2848
rect 437523 2808 476212 2836
rect 437523 2805 437535 2808
rect 437477 2799 437535 2805
rect 476206 2796 476212 2808
rect 476264 2796 476270 2848
rect 502058 2796 502064 2848
rect 502116 2836 502122 2848
rect 529014 2836 529020 2848
rect 502116 2808 529020 2836
rect 502116 2796 502122 2808
rect 529014 2796 529020 2808
rect 529072 2796 529078 2848
rect 1104 2672 582820 2768
rect 126885 2635 126943 2641
rect 126885 2601 126897 2635
rect 126931 2632 126943 2635
rect 132313 2635 132371 2641
rect 132313 2632 132325 2635
rect 126931 2604 132325 2632
rect 126931 2601 126943 2604
rect 126885 2595 126943 2601
rect 132313 2601 132325 2604
rect 132359 2601 132371 2635
rect 132313 2595 132371 2601
rect 440326 2592 440332 2644
rect 440384 2632 440390 2644
rect 441706 2632 441712 2644
rect 440384 2604 441712 2632
rect 440384 2592 440390 2604
rect 441706 2592 441712 2604
rect 441764 2592 441770 2644
rect 447410 2592 447416 2644
rect 447468 2632 447474 2644
rect 460753 2635 460811 2641
rect 460753 2632 460765 2635
rect 447468 2604 460765 2632
rect 447468 2592 447474 2604
rect 460753 2601 460765 2604
rect 460799 2601 460811 2635
rect 460753 2595 460811 2601
rect 518897 2635 518955 2641
rect 518897 2601 518909 2635
rect 518943 2632 518955 2635
rect 525426 2632 525432 2644
rect 518943 2604 525432 2632
rect 518943 2601 518955 2604
rect 518897 2595 518955 2601
rect 525426 2592 525432 2604
rect 525484 2592 525490 2644
rect 121086 2524 121092 2576
rect 121144 2564 121150 2576
rect 128449 2567 128507 2573
rect 128449 2564 128461 2567
rect 121144 2536 128461 2564
rect 121144 2524 121150 2536
rect 128449 2533 128461 2536
rect 128495 2533 128507 2567
rect 128449 2527 128507 2533
rect 1104 2128 582820 2224
rect 340874 1980 340880 2032
rect 340932 2020 340938 2032
rect 342162 2020 342168 2032
rect 340932 1992 342168 2020
rect 340932 1980 340938 1992
rect 342162 1980 342168 1992
rect 342220 1980 342226 2032
<< via1 >>
rect 40500 700476 40552 700528
rect 41328 700476 41380 700528
rect 480168 700476 480220 700528
rect 527180 700476 527232 700528
rect 402888 700408 402940 700460
rect 429844 700408 429896 700460
rect 441528 700408 441580 700460
rect 478512 700408 478564 700460
rect 492588 700408 492640 700460
rect 543464 700408 543516 700460
rect 378048 700340 378100 700392
rect 397460 700340 397512 700392
rect 416688 700340 416740 700392
rect 446128 700340 446180 700392
rect 453948 700340 454000 700392
rect 494796 700340 494848 700392
rect 506388 700340 506440 700392
rect 559656 700340 559708 700392
rect 56784 700272 56836 700324
rect 57888 700272 57940 700324
rect 186504 700272 186556 700324
rect 187608 700272 187660 700324
rect 339408 700272 339460 700324
rect 348792 700272 348844 700324
rect 351828 700272 351880 700324
rect 364984 700272 365036 700324
rect 365628 700272 365680 700324
rect 381176 700272 381228 700324
rect 390468 700272 390520 700324
rect 413652 700272 413704 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 467748 700272 467800 700324
rect 510988 700272 511040 700324
rect 517428 700272 517480 700324
rect 575848 700272 575900 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 251456 699660 251508 699712
rect 252468 699660 252520 699712
rect 299480 699660 299532 699712
rect 300124 699660 300176 699712
rect 313188 699660 313240 699712
rect 316316 699660 316368 699712
rect 326988 699660 327040 699712
rect 332508 699660 332560 699712
rect 520924 696940 520976 696992
rect 580172 696940 580224 696992
rect 521016 683136 521068 683188
rect 580172 683136 580224 683188
rect 284208 682864 284260 682916
rect 287612 682864 287664 682916
rect 57888 682592 57940 682644
rect 108396 682592 108448 682644
rect 41328 682524 41380 682576
rect 95608 682524 95660 682576
rect 106188 682524 106240 682576
rect 146852 682524 146904 682576
rect 154488 682524 154540 682576
rect 185216 682524 185268 682576
rect 24768 682456 24820 682508
rect 82820 682456 82872 682508
rect 89628 682456 89680 682508
rect 134064 682456 134116 682508
rect 137928 682456 137980 682508
rect 172428 682456 172480 682508
rect 187608 682456 187660 682508
rect 210792 682456 210844 682508
rect 219348 682456 219400 682508
rect 236368 682456 236420 682508
rect 8208 682388 8260 682440
rect 71044 682388 71096 682440
rect 73068 682388 73120 682440
rect 121184 682388 121236 682440
rect 122748 682388 122800 682440
rect 159640 682388 159692 682440
rect 171048 682388 171100 682440
rect 198004 682388 198056 682440
rect 202788 682388 202840 682440
rect 223580 682388 223632 682440
rect 235908 682388 235960 682440
rect 249248 682388 249300 682440
rect 252468 682388 252520 682440
rect 262036 682388 262088 682440
rect 267648 682388 267700 682440
rect 274824 682388 274876 682440
rect 325976 681708 326028 681760
rect 326988 681708 327040 681760
rect 338764 681708 338816 681760
rect 339408 681708 339460 681760
rect 364432 681708 364484 681760
rect 365628 681708 365680 681760
rect 377220 681708 377272 681760
rect 378048 681708 378100 681760
rect 390008 681708 390060 681760
rect 390468 681708 390520 681760
rect 415584 681708 415636 681760
rect 416688 681708 416740 681760
rect 428372 681708 428424 681760
rect 429108 681708 429160 681760
rect 466736 681708 466788 681760
rect 467748 681708 467800 681760
rect 479616 681708 479668 681760
rect 480168 681708 480220 681760
rect 505192 681708 505244 681760
rect 506388 681708 506440 681760
rect 3424 680280 3476 680332
rect 66996 680280 67048 680332
rect 520924 670828 520976 670880
rect 580172 670828 580224 670880
rect 3516 669264 3568 669316
rect 67180 669264 67232 669316
rect 3424 658112 3476 658164
rect 67364 658112 67416 658164
rect 521016 656888 521068 656940
rect 580172 656888 580224 656940
rect 3516 647164 3568 647216
rect 67364 647164 67416 647216
rect 520924 643084 520976 643136
rect 580172 643084 580224 643136
rect 3424 636148 3476 636200
rect 67364 636148 67416 636200
rect 520924 630640 520976 630692
rect 580172 630640 580224 630692
rect 3424 624928 3476 624980
rect 67364 624928 67416 624980
rect 520280 616972 520332 617024
rect 580172 616972 580224 617024
rect 3424 614048 3476 614100
rect 66904 614048 66956 614100
rect 521108 603100 521160 603152
rect 580172 603100 580224 603152
rect 4068 603032 4120 603084
rect 66444 603032 66496 603084
rect 3424 591948 3476 592000
rect 66996 591948 67048 592000
rect 521568 590656 521620 590708
rect 579804 590656 579856 590708
rect 3424 579572 3476 579624
rect 67180 579572 67232 579624
rect 521568 577464 521620 577516
rect 580172 577464 580224 577516
rect 4068 567196 4120 567248
rect 67364 567196 67416 567248
rect 520740 564340 520792 564392
rect 580172 564340 580224 564392
rect 3424 556180 3476 556232
rect 67364 556180 67416 556232
rect 521016 551964 521068 552016
rect 579988 551964 580040 552016
rect 2964 545164 3016 545216
rect 66628 545164 66680 545216
rect 520924 538160 520976 538212
rect 580172 538160 580224 538212
rect 3424 534080 3476 534132
rect 67364 534080 67416 534132
rect 520924 525716 520976 525768
rect 579804 525716 579856 525768
rect 3424 522996 3476 523048
rect 66444 522996 66496 523048
rect 3424 511980 3476 512032
rect 67364 511980 67416 512032
rect 520924 511776 520976 511828
rect 580172 511776 580224 511828
rect 3516 501100 3568 501152
rect 67456 501100 67508 501152
rect 521016 498108 521068 498160
rect 580172 498108 580224 498160
rect 3424 489880 3476 489932
rect 67456 489880 67508 489932
rect 520924 485664 520976 485716
rect 580172 485664 580224 485716
rect 3516 478864 3568 478916
rect 67364 478864 67416 478916
rect 521016 471928 521068 471980
rect 580172 471928 580224 471980
rect 3424 466420 3476 466472
rect 66996 466420 67048 466472
rect 520924 458124 520976 458176
rect 580172 458124 580224 458176
rect 3516 455404 3568 455456
rect 67364 455404 67416 455456
rect 521108 445680 521160 445732
rect 580172 445680 580224 445732
rect 3424 444524 3476 444576
rect 66720 444524 66772 444576
rect 3608 433304 3660 433356
rect 67180 433304 67232 433356
rect 521016 431808 521068 431860
rect 580172 431808 580224 431860
rect 3516 422288 3568 422340
rect 66812 422288 66864 422340
rect 520924 419296 520976 419348
rect 580172 419296 580224 419348
rect 3424 411340 3476 411392
rect 67272 411340 67324 411392
rect 521016 405628 521068 405680
rect 580172 405628 580224 405680
rect 3608 400188 3660 400240
rect 67456 400188 67508 400240
rect 520924 391892 520976 391944
rect 580172 391892 580224 391944
rect 3516 389172 3568 389224
rect 67364 389172 67416 389224
rect 521108 379448 521160 379500
rect 580172 379448 580224 379500
rect 3424 378156 3476 378208
rect 67364 378156 67416 378208
rect 3700 367072 3752 367124
rect 67364 367072 67416 367124
rect 521016 365644 521068 365696
rect 580172 365644 580224 365696
rect 3608 356056 3660 356108
rect 67364 356056 67416 356108
rect 520924 353200 520976 353252
rect 580172 353200 580224 353252
rect 3516 343612 3568 343664
rect 67364 343612 67416 343664
rect 521200 339328 521252 339380
rect 580172 339328 580224 339380
rect 3424 332596 3476 332648
rect 67180 332596 67232 332648
rect 521108 325592 521160 325644
rect 580172 325592 580224 325644
rect 3700 321580 3752 321632
rect 67364 321580 67416 321632
rect 521016 313216 521068 313268
rect 580172 313216 580224 313268
rect 3608 310496 3660 310548
rect 66720 310496 66772 310548
rect 3516 299480 3568 299532
rect 67364 299480 67416 299532
rect 520924 299412 520976 299464
rect 580172 299412 580224 299464
rect 3424 288396 3476 288448
rect 66444 288396 66496 288448
rect 521200 285472 521252 285524
rect 580172 285472 580224 285524
rect 3792 277516 3844 277568
rect 67364 277516 67416 277568
rect 521108 273164 521160 273216
rect 580172 273164 580224 273216
rect 3700 266364 3752 266416
rect 67364 266364 67416 266416
rect 521016 259360 521068 259412
rect 580172 259360 580224 259412
rect 3608 255280 3660 255332
rect 67364 255280 67416 255332
rect 520924 245556 520976 245608
rect 580172 245556 580224 245608
rect 3516 244332 3568 244384
rect 67364 244332 67416 244384
rect 3424 233248 3476 233300
rect 67180 233248 67232 233300
rect 521292 233180 521344 233232
rect 579988 233180 580040 233232
rect 3884 220940 3936 220992
rect 67364 220940 67416 220992
rect 521200 219376 521252 219428
rect 580172 219376 580224 219428
rect 3792 209788 3844 209840
rect 67364 209788 67416 209840
rect 521108 206932 521160 206984
rect 579804 206932 579856 206984
rect 3700 198704 3752 198756
rect 67364 198704 67416 198756
rect 521016 192992 521068 193044
rect 580172 192992 580224 193044
rect 3608 187756 3660 187808
rect 67456 187756 67508 187808
rect 520924 179324 520976 179376
rect 580172 179324 580224 179376
rect 3516 176672 3568 176724
rect 67364 176672 67416 176724
rect 521384 166880 521436 166932
rect 580172 166880 580224 166932
rect 3424 165588 3476 165640
rect 67364 165588 67416 165640
rect 3976 154572 4028 154624
rect 67272 154572 67324 154624
rect 521292 153144 521344 153196
rect 580172 153144 580224 153196
rect 3884 143692 3936 143744
rect 67364 143692 67416 143744
rect 521200 139340 521252 139392
rect 580172 139340 580224 139392
rect 3792 132472 3844 132524
rect 67180 132472 67232 132524
rect 521108 126896 521160 126948
rect 580172 126896 580224 126948
rect 3700 121456 3752 121508
rect 67364 121456 67416 121508
rect 521016 113024 521068 113076
rect 580172 113024 580224 113076
rect 3608 109012 3660 109064
rect 67364 109012 67416 109064
rect 520924 100512 520976 100564
rect 580172 100512 580224 100564
rect 3516 97996 3568 98048
rect 67180 97996 67232 98048
rect 3424 88340 3476 88392
rect 67456 88340 67508 88392
rect 73160 87796 73212 87848
rect 74436 87796 74488 87848
rect 78680 87796 78732 87848
rect 79956 87796 80008 87848
rect 110420 87796 110472 87848
rect 111696 87796 111748 87848
rect 116032 87796 116084 87848
rect 117216 87796 117268 87848
rect 147772 87796 147824 87848
rect 148956 87796 149008 87848
rect 150532 87796 150584 87848
rect 151716 87796 151768 87848
rect 158720 87796 158772 87848
rect 159904 87796 159956 87848
rect 167000 87796 167052 87848
rect 168092 87796 168144 87848
rect 169760 87796 169812 87848
rect 170760 87796 170812 87848
rect 296720 87796 296772 87848
rect 297996 87796 298048 87848
rect 299480 87796 299532 87848
rect 300756 87796 300808 87848
rect 316040 87796 316092 87848
rect 317040 87796 317092 87848
rect 321560 87796 321612 87848
rect 322560 87796 322612 87848
rect 333980 87796 334032 87848
rect 335256 87796 335308 87848
rect 402980 87796 403032 87848
rect 404256 87796 404308 87848
rect 405740 87796 405792 87848
rect 407016 87796 407068 87848
rect 408500 87796 408552 87848
rect 409776 87796 409828 87848
rect 422300 87796 422352 87848
rect 423392 87796 423444 87848
rect 430580 87796 430632 87848
rect 431580 87796 431632 87848
rect 443092 87796 443144 87848
rect 444276 87796 444328 87848
rect 448520 87796 448572 87848
rect 449704 87796 449756 87848
rect 454040 87796 454092 87848
rect 455132 87796 455184 87848
rect 456800 87796 456852 87848
rect 457892 87796 457944 87848
rect 459652 87796 459704 87848
rect 460652 87796 460704 87848
rect 521476 86912 521528 86964
rect 580172 86912 580224 86964
rect 76012 86096 76064 86148
rect 77208 86096 77260 86148
rect 103520 86096 103572 86148
rect 104440 86096 104492 86148
rect 106280 86096 106332 86148
rect 107200 86096 107252 86148
rect 109040 86096 109092 86148
rect 109960 86096 110012 86148
rect 140780 86096 140832 86148
rect 141700 86096 141752 86148
rect 294052 86096 294104 86148
rect 295248 86096 295300 86148
rect 331312 86096 331364 86148
rect 332508 86096 332560 86148
rect 438860 86096 438912 86148
rect 439780 86096 439832 86148
rect 445852 86096 445904 86148
rect 447048 86096 447100 86148
rect 76564 85484 76616 85536
rect 78128 85484 78180 85536
rect 79324 85484 79376 85536
rect 80888 85484 80940 85536
rect 94504 85484 94556 85536
rect 95148 85484 95200 85536
rect 95424 85484 95476 85536
rect 96436 85484 96488 85536
rect 97172 85484 97224 85536
rect 97908 85484 97960 85536
rect 98092 85484 98144 85536
rect 99288 85484 99340 85536
rect 99932 85484 99984 85536
rect 100668 85484 100720 85536
rect 100852 85484 100904 85536
rect 102048 85484 102100 85536
rect 115204 85484 115256 85536
rect 116308 85484 116360 85536
rect 119344 85484 119396 85536
rect 120816 85484 120868 85536
rect 130384 85484 130436 85536
rect 131764 85484 131816 85536
rect 146944 85484 146996 85536
rect 148048 85484 148100 85536
rect 176016 85484 176068 85536
rect 177120 85484 177172 85536
rect 180800 85484 180852 85536
rect 182180 85484 182232 85536
rect 182640 85484 182692 85536
rect 184204 85484 184256 85536
rect 184388 85484 184440 85536
rect 186964 85484 187016 85536
rect 187148 85484 187200 85536
rect 187608 85484 187660 85536
rect 188068 85484 188120 85536
rect 188988 85484 189040 85536
rect 190828 85484 190880 85536
rect 191656 85484 191708 85536
rect 192576 85484 192628 85536
rect 193128 85484 193180 85536
rect 193496 85484 193548 85536
rect 194508 85484 194560 85536
rect 195336 85484 195388 85536
rect 195888 85484 195940 85536
rect 196256 85484 196308 85536
rect 197176 85484 197228 85536
rect 198096 85484 198148 85536
rect 198648 85484 198700 85536
rect 198924 85484 198976 85536
rect 199936 85484 199988 85536
rect 200764 85484 200816 85536
rect 201408 85484 201460 85536
rect 201684 85484 201736 85536
rect 202788 85484 202840 85536
rect 203524 85484 203576 85536
rect 204168 85484 204220 85536
rect 204444 85484 204496 85536
rect 205456 85484 205508 85536
rect 206192 85484 206244 85536
rect 206928 85484 206980 85536
rect 208952 85484 209004 85536
rect 209688 85484 209740 85536
rect 211712 85484 211764 85536
rect 212448 85484 212500 85536
rect 212632 85484 212684 85536
rect 213828 85484 213880 85536
rect 214380 85484 214432 85536
rect 215208 85484 215260 85536
rect 215300 85484 215352 85536
rect 216588 85484 216640 85536
rect 217140 85484 217192 85536
rect 217968 85484 218020 85536
rect 218060 85484 218112 85536
rect 219348 85484 219400 85536
rect 219900 85484 219952 85536
rect 220728 85484 220780 85536
rect 222568 85484 222620 85536
rect 223488 85484 223540 85536
rect 224408 85484 224460 85536
rect 224868 85484 224920 85536
rect 225328 85484 225380 85536
rect 226156 85484 226208 85536
rect 227168 85484 227220 85536
rect 227628 85484 227680 85536
rect 229836 85484 229888 85536
rect 230296 85484 230348 85536
rect 230756 85484 230808 85536
rect 231768 85484 231820 85536
rect 232596 85484 232648 85536
rect 233148 85484 233200 85536
rect 233516 85484 233568 85536
rect 234436 85484 234488 85536
rect 235264 85484 235316 85536
rect 235908 85484 235960 85536
rect 236184 85484 236236 85536
rect 237196 85484 237248 85536
rect 238024 85484 238076 85536
rect 238668 85484 238720 85536
rect 240784 85484 240836 85536
rect 241336 85484 241388 85536
rect 241704 85484 241756 85536
rect 242716 85484 242768 85536
rect 243452 85484 243504 85536
rect 244188 85484 244240 85536
rect 244372 85484 244424 85536
rect 245568 85484 245620 85536
rect 246212 85484 246264 85536
rect 246948 85484 247000 85536
rect 247132 85484 247184 85536
rect 248328 85484 248380 85536
rect 248972 85484 249024 85536
rect 249708 85484 249760 85536
rect 249800 85484 249852 85536
rect 251088 85484 251140 85536
rect 251640 85484 251692 85536
rect 252468 85484 252520 85536
rect 252560 85484 252612 85536
rect 253848 85484 253900 85536
rect 254400 85484 254452 85536
rect 255228 85484 255280 85536
rect 255320 85484 255372 85536
rect 256608 85484 256660 85536
rect 256700 85484 256752 85536
rect 257988 85484 258040 85536
rect 258080 85484 258132 85536
rect 258908 85484 258960 85536
rect 259828 85484 259880 85536
rect 260748 85484 260800 85536
rect 262588 85484 262640 85536
rect 263508 85484 263560 85536
rect 264336 85484 264388 85536
rect 264888 85484 264940 85536
rect 265256 85484 265308 85536
rect 266268 85484 266320 85536
rect 267096 85484 267148 85536
rect 267648 85484 267700 85536
rect 268016 85484 268068 85536
rect 269028 85484 269080 85536
rect 269856 85484 269908 85536
rect 270408 85484 270460 85536
rect 270776 85484 270828 85536
rect 271788 85484 271840 85536
rect 272524 85484 272576 85536
rect 273168 85484 273220 85536
rect 273444 85484 273496 85536
rect 274548 85484 274600 85536
rect 275284 85484 275336 85536
rect 275928 85484 275980 85536
rect 276204 85484 276256 85536
rect 277216 85484 277268 85536
rect 278044 85484 278096 85536
rect 278688 85484 278740 85536
rect 278964 85484 279016 85536
rect 280068 85484 280120 85536
rect 280160 85484 280212 85536
rect 280712 85484 280764 85536
rect 280804 85484 280856 85536
rect 282552 85484 282604 85536
rect 289084 85484 289136 85536
rect 289820 85484 289872 85536
rect 308404 85484 308456 85536
rect 309784 85484 309836 85536
rect 309876 85484 309928 85536
rect 310704 85484 310756 85536
rect 312544 85484 312596 85536
rect 313464 85484 313516 85536
rect 337108 85484 337160 85536
rect 338028 85484 338080 85536
rect 338856 85484 338908 85536
rect 339408 85484 339460 85536
rect 339776 85484 339828 85536
rect 340788 85484 340840 85536
rect 341616 85484 341668 85536
rect 342168 85484 342220 85536
rect 342536 85484 342588 85536
rect 343456 85484 343508 85536
rect 344376 85484 344428 85536
rect 344928 85484 344980 85536
rect 345204 85484 345256 85536
rect 346308 85484 346360 85536
rect 347044 85484 347096 85536
rect 347688 85484 347740 85536
rect 347964 85484 348016 85536
rect 348976 85484 349028 85536
rect 349804 85484 349856 85536
rect 350448 85484 350500 85536
rect 350724 85484 350776 85536
rect 351828 85484 351880 85536
rect 353392 85484 353444 85536
rect 354496 85484 354548 85536
rect 355232 85484 355284 85536
rect 355968 85484 356020 85536
rect 356152 85484 356204 85536
rect 357256 85484 357308 85536
rect 357992 85484 358044 85536
rect 358728 85484 358780 85536
rect 358912 85484 358964 85536
rect 360016 85484 360068 85536
rect 360660 85484 360712 85536
rect 361488 85484 361540 85536
rect 361580 85484 361632 85536
rect 362868 85484 362920 85536
rect 363420 85484 363472 85536
rect 364248 85484 364300 85536
rect 364340 85484 364392 85536
rect 365536 85484 365588 85536
rect 366180 85484 366232 85536
rect 367008 85484 367060 85536
rect 367928 85484 367980 85536
rect 368388 85484 368440 85536
rect 368848 85484 368900 85536
rect 369768 85484 369820 85536
rect 370688 85484 370740 85536
rect 371148 85484 371200 85536
rect 371608 85484 371660 85536
rect 372436 85484 372488 85536
rect 374276 85484 374328 85536
rect 375196 85484 375248 85536
rect 376116 85484 376168 85536
rect 376668 85484 376720 85536
rect 377036 85484 377088 85536
rect 378048 85484 378100 85536
rect 378876 85484 378928 85536
rect 379428 85484 379480 85536
rect 379796 85484 379848 85536
rect 380808 85484 380860 85536
rect 381636 85484 381688 85536
rect 382188 85484 382240 85536
rect 382464 85484 382516 85536
rect 383476 85484 383528 85536
rect 384304 85484 384356 85536
rect 384948 85484 385000 85536
rect 385224 85484 385276 85536
rect 386236 85484 386288 85536
rect 387064 85484 387116 85536
rect 387708 85484 387760 85536
rect 387984 85484 388036 85536
rect 389088 85484 389140 85536
rect 389732 85484 389784 85536
rect 390468 85484 390520 85536
rect 390652 85484 390704 85536
rect 391848 85484 391900 85536
rect 392492 85484 392544 85536
rect 393228 85484 393280 85536
rect 393412 85484 393464 85536
rect 394608 85484 394660 85536
rect 395252 85484 395304 85536
rect 395988 85484 396040 85536
rect 396172 85484 396224 85536
rect 397276 85484 397328 85536
rect 397920 85484 397972 85536
rect 398748 85484 398800 85536
rect 401508 85484 401560 85536
rect 402520 85484 402572 85536
rect 435364 85484 435416 85536
rect 436100 85484 436152 85536
rect 439504 85484 439556 85536
rect 441528 85484 441580 85536
rect 442264 85484 442316 85536
rect 443368 85484 443420 85536
rect 462228 85484 462280 85536
rect 484308 85484 484360 85536
rect 493324 85484 493376 85536
rect 493968 85484 494020 85536
rect 494244 85484 494296 85536
rect 495348 85484 495400 85536
rect 496084 85484 496136 85536
rect 496728 85484 496780 85536
rect 497004 85484 497056 85536
rect 498108 85484 498160 85536
rect 498844 85484 498896 85536
rect 499488 85484 499540 85536
rect 499672 85484 499724 85536
rect 500776 85484 500828 85536
rect 501512 85484 501564 85536
rect 502248 85484 502300 85536
rect 502432 85484 502484 85536
rect 503536 85484 503588 85536
rect 504272 85484 504324 85536
rect 505008 85484 505060 85536
rect 505192 85484 505244 85536
rect 506296 85484 506348 85536
rect 506940 85484 506992 85536
rect 507768 85484 507820 85536
rect 507860 85484 507912 85536
rect 509056 85484 509108 85536
rect 509700 85484 509752 85536
rect 510528 85484 510580 85536
rect 510620 85484 510672 85536
rect 511816 85484 511868 85536
rect 512460 85484 512512 85536
rect 513288 85484 513340 85536
rect 514208 85484 514260 85536
rect 514668 85484 514720 85536
rect 515128 85484 515180 85536
rect 516048 85484 516100 85536
rect 516968 85484 517020 85536
rect 517428 85484 517480 85536
rect 517888 85484 517940 85536
rect 518808 85484 518860 85536
rect 175924 85280 175976 85332
rect 178040 85280 178092 85332
rect 183560 85280 183612 85332
rect 184848 85280 184900 85332
rect 207112 85280 207164 85332
rect 209044 85280 209096 85332
rect 209872 85280 209924 85332
rect 214564 85280 214616 85332
rect 221648 85280 221700 85332
rect 224224 85280 224276 85332
rect 238944 85280 238996 85332
rect 240784 85280 240836 85332
rect 261668 85280 261720 85332
rect 267004 85280 267056 85332
rect 279792 85280 279844 85332
rect 280896 85280 280948 85332
rect 281632 85280 281684 85332
rect 286416 85280 286468 85332
rect 310428 85280 310480 85332
rect 311624 85280 311676 85332
rect 351644 85280 351696 85332
rect 352656 85280 352708 85332
rect 455328 85280 455380 85332
rect 482468 85280 482520 85332
rect 482928 85280 482980 85332
rect 489736 85280 489788 85332
rect 513380 85280 513432 85332
rect 514576 85280 514628 85332
rect 107568 85212 107620 85264
rect 155316 85212 155368 85264
rect 451188 85212 451240 85264
rect 481548 85212 481600 85264
rect 96528 85144 96580 85196
rect 152648 85144 152700 85196
rect 161388 85144 161440 85196
rect 175372 85144 175424 85196
rect 444288 85144 444340 85196
rect 479708 85144 479760 85196
rect 18604 85076 18656 85128
rect 132592 85076 132644 85128
rect 151728 85076 151780 85128
rect 172612 85076 172664 85128
rect 437388 85076 437440 85128
rect 477868 85076 477920 85128
rect 480168 85076 480220 85128
rect 488816 85076 488868 85128
rect 19984 85008 20036 85060
rect 161664 85008 161716 85060
rect 352472 85008 352524 85060
rect 398104 85008 398156 85060
rect 423588 85008 423640 85060
rect 474280 85008 474332 85060
rect 476028 85008 476080 85060
rect 487896 85008 487948 85060
rect 7564 84940 7616 84992
rect 165344 84940 165396 84992
rect 165528 84940 165580 84992
rect 176292 84940 176344 84992
rect 189908 84940 189960 84992
rect 195244 84940 195296 84992
rect 228916 84940 228968 84992
rect 232504 84940 232556 84992
rect 239864 84940 239916 84992
rect 249064 84940 249116 84992
rect 254584 84940 254636 84992
rect 286232 84940 286284 84992
rect 287704 84940 287756 84992
rect 401600 84940 401652 84992
rect 416688 84940 416740 84992
rect 472440 84940 472492 84992
rect 473268 84940 473320 84992
rect 486976 84940 487028 84992
rect 495164 84940 495216 84992
rect 503812 84940 503864 84992
rect 466368 84736 466420 84788
rect 485136 84736 485188 84788
rect 469128 84668 469180 84720
rect 486056 84668 486108 84720
rect 227996 84600 228048 84652
rect 229744 84600 229796 84652
rect 373448 84600 373500 84652
rect 376024 84600 376076 84652
rect 208032 84396 208084 84448
rect 211804 84396 211856 84448
rect 112444 84192 112496 84244
rect 114468 84192 114520 84244
rect 169024 84192 169076 84244
rect 171692 84192 171744 84244
rect 257068 84192 257120 84244
rect 258724 84192 258776 84244
rect 286324 84192 286376 84244
rect 287060 84192 287112 84244
rect 487068 84192 487120 84244
rect 490656 84192 490708 84244
rect 62028 83512 62080 83564
rect 84292 83512 84344 83564
rect 153108 83512 153160 83564
rect 288440 83512 288492 83564
rect 292488 83512 292540 83564
rect 440332 83512 440384 83564
rect 10324 83444 10376 83496
rect 71872 83444 71924 83496
rect 129648 83444 129700 83496
rect 167092 83444 167144 83496
rect 184940 83444 184992 83496
rect 200120 83444 200172 83496
rect 256700 83444 256752 83496
rect 483112 83444 483164 83496
rect 309784 82220 309836 82272
rect 444380 82220 444432 82272
rect 241428 80792 241480 80844
rect 310428 80792 310480 80844
rect 59268 80724 59320 80776
rect 84108 80724 84160 80776
rect 133788 80724 133840 80776
rect 167000 80724 167052 80776
rect 258080 80724 258132 80776
rect 487160 80724 487212 80776
rect 14464 80656 14516 80708
rect 102140 80656 102192 80708
rect 143448 80656 143500 80708
rect 401508 80656 401560 80708
rect 344836 79296 344888 79348
rect 454132 79296 454184 79348
rect 230388 78072 230440 78124
rect 307852 78072 307904 78124
rect 70216 78004 70268 78056
rect 116032 78004 116084 78056
rect 137928 78004 137980 78056
rect 284392 78004 284444 78056
rect 352564 78004 352616 78056
rect 455420 78004 455472 78056
rect 12348 77936 12400 77988
rect 73252 77936 73304 77988
rect 280160 77936 280212 77988
rect 572720 77936 572772 77988
rect 281448 76508 281500 76560
rect 437480 76508 437532 76560
rect 227536 75284 227588 75336
rect 307760 75284 307812 75336
rect 30288 75216 30340 75268
rect 76012 75216 76064 75268
rect 155868 75216 155920 75268
rect 289084 75216 289136 75268
rect 75828 75148 75880 75200
rect 146392 75148 146444 75200
rect 280896 75148 280948 75200
rect 568580 75148 568632 75200
rect 224224 74060 224276 74112
rect 340880 74060 340932 74112
rect 148968 73856 149020 73908
rect 287152 73856 287204 73908
rect 375196 73856 375248 73908
rect 484400 73856 484452 73908
rect 34428 73788 34480 73840
rect 76564 73788 76616 73840
rect 92388 73788 92440 73840
rect 121552 73788 121604 73840
rect 274364 73788 274416 73840
rect 435364 73788 435416 73840
rect 521384 73108 521436 73160
rect 580172 73108 580224 73160
rect 220636 71068 220688 71120
rect 338120 71068 338172 71120
rect 37188 71000 37240 71052
rect 78772 71000 78824 71052
rect 255228 71000 255280 71052
rect 469312 71000 469364 71052
rect 220728 68348 220780 68400
rect 334164 68348 334216 68400
rect 15844 68280 15896 68332
rect 103612 68280 103664 68332
rect 253756 68280 253808 68332
rect 465264 68280 465316 68332
rect 252284 66988 252336 67040
rect 430672 66988 430724 67040
rect 219256 65560 219308 65612
rect 331404 65560 331456 65612
rect 349804 65560 349856 65612
rect 454040 65560 454092 65612
rect 28908 65492 28960 65544
rect 106372 65492 106424 65544
rect 252468 65492 252520 65544
rect 458272 65492 458324 65544
rect 358084 64268 358136 64320
rect 456892 64268 456944 64320
rect 219348 62908 219400 62960
rect 327264 62908 327316 62960
rect 324228 62840 324280 62892
rect 448612 62840 448664 62892
rect 32404 62772 32456 62824
rect 106280 62772 106332 62824
rect 241336 62772 241388 62824
rect 415492 62772 415544 62824
rect 146208 61344 146260 61396
rect 403072 61344 403124 61396
rect 521292 60664 521344 60716
rect 580172 60664 580224 60716
rect 217968 60120 218020 60172
rect 324504 60120 324556 60172
rect 318064 60052 318116 60104
rect 445852 60052 445904 60104
rect 38568 59984 38620 60036
rect 109132 59984 109184 60036
rect 249064 59984 249116 60036
rect 412732 59984 412784 60036
rect 278044 58624 278096 58676
rect 436192 58624 436244 58676
rect 216496 57332 216548 57384
rect 320272 57332 320324 57384
rect 308496 57264 308548 57316
rect 443092 57264 443144 57316
rect 10968 57196 11020 57248
rect 130384 57196 130436 57248
rect 238668 57196 238720 57248
rect 405924 57196 405976 57248
rect 216588 56108 216640 56160
rect 316224 56108 316276 56160
rect 299388 55904 299440 55956
rect 441620 55904 441672 55956
rect 50988 55836 51040 55888
rect 140872 55836 140924 55888
rect 237196 55836 237248 55888
rect 399024 55836 399076 55888
rect 235816 54476 235868 54528
rect 425152 54476 425204 54528
rect 215208 53184 215260 53236
rect 313372 53184 313424 53236
rect 285588 53116 285640 53168
rect 438952 53116 439004 53168
rect 57888 53048 57940 53100
rect 142160 53048 142212 53100
rect 235908 53048 235960 53100
rect 394700 53048 394752 53100
rect 267556 51756 267608 51808
rect 433432 51756 433484 51808
rect 213736 50396 213788 50448
rect 309140 50396 309192 50448
rect 377956 50396 378008 50448
rect 485044 50396 485096 50448
rect 64788 50328 64840 50380
rect 143632 50328 143684 50380
rect 234436 50328 234488 50380
rect 387800 50328 387852 50380
rect 263324 49036 263376 49088
rect 433340 49036 433392 49088
rect 213828 47608 213880 47660
rect 306472 47608 306524 47660
rect 378048 47608 378100 47660
rect 487804 47608 487856 47660
rect 61936 47540 61988 47592
rect 143540 47540 143592 47592
rect 233148 47540 233200 47592
rect 383660 47540 383712 47592
rect 521200 46860 521252 46912
rect 580172 46860 580224 46912
rect 256424 46316 256476 46368
rect 430580 46316 430632 46368
rect 344284 44956 344336 45008
rect 452660 44956 452712 45008
rect 212448 44888 212500 44940
rect 302424 44888 302476 44940
rect 376668 44888 376720 44940
rect 489184 44888 489236 44940
rect 68928 44820 68980 44872
rect 144920 44820 144972 44872
rect 231676 44820 231728 44872
rect 380900 44820 380952 44872
rect 231676 43392 231728 43444
rect 425060 43392 425112 43444
rect 338764 42168 338816 42220
rect 451372 42168 451424 42220
rect 211068 42100 211120 42152
rect 299664 42100 299716 42152
rect 375288 42100 375340 42152
rect 488540 42100 488592 42152
rect 53748 42032 53800 42084
rect 140780 42032 140832 42084
rect 231768 42032 231820 42084
rect 376760 42032 376812 42084
rect 249616 40672 249668 40724
rect 429200 40672 429252 40724
rect 214564 39380 214616 39432
rect 295432 39380 295484 39432
rect 336004 39380 336056 39432
rect 451280 39380 451332 39432
rect 71688 39312 71740 39364
rect 146300 39312 146352 39364
rect 230296 39312 230348 39364
rect 374000 39312 374052 39364
rect 376024 39312 376076 39364
rect 481640 39312 481692 39364
rect 211804 38156 211856 38208
rect 288440 38156 288492 38208
rect 232504 37952 232556 38004
rect 369860 37952 369912 38004
rect 35808 37884 35860 37936
rect 107660 37884 107712 37936
rect 256516 37884 256568 37936
rect 476304 37884 476356 37936
rect 245384 36524 245436 36576
rect 427912 36524 427964 36576
rect 209044 35436 209096 35488
rect 284484 35436 284536 35488
rect 288348 35232 288400 35284
rect 438860 35232 438912 35284
rect 45468 35164 45520 35216
rect 110512 35164 110564 35216
rect 135168 35164 135220 35216
rect 284300 35164 284352 35216
rect 286416 35164 286468 35216
rect 575480 35164 575532 35216
rect 242624 33804 242676 33856
rect 427820 33804 427872 33856
rect 521108 33056 521160 33108
rect 580172 33056 580224 33108
rect 206928 32512 206980 32564
rect 281540 32512 281592 32564
rect 229744 32444 229796 32496
rect 365720 32444 365772 32496
rect 23388 32376 23440 32428
rect 104900 32376 104952 32428
rect 117228 32376 117280 32428
rect 128360 32376 128412 32428
rect 256608 32376 256660 32428
rect 473452 32376 473504 32428
rect 237196 31084 237248 31136
rect 309876 31084 309928 31136
rect 331128 31084 331180 31136
rect 449900 31084 449952 31136
rect 223304 29724 223356 29776
rect 306380 29724 306432 29776
rect 144828 29656 144880 29708
rect 286324 29656 286376 29708
rect 326988 29656 327040 29708
rect 448520 29656 448572 29708
rect 19248 29588 19300 29640
rect 103520 29588 103572 29640
rect 113088 29588 113140 29640
rect 127072 29588 127124 29640
rect 264888 29588 264940 29640
rect 507860 29588 507912 29640
rect 248144 28364 248196 28416
rect 312544 28364 312596 28416
rect 320824 28364 320876 28416
rect 447140 28364 447192 28416
rect 95056 26936 95108 26988
rect 122840 26936 122892 26988
rect 162768 26936 162820 26988
rect 291200 26936 291252 26988
rect 295248 26936 295300 26988
rect 439504 26936 439556 26988
rect 42708 26868 42760 26920
rect 109040 26868 109092 26920
rect 263416 26868 263468 26920
rect 505100 26868 505152 26920
rect 124128 26460 124180 26512
rect 129832 26460 129884 26512
rect 244096 25644 244148 25696
rect 311900 25644 311952 25696
rect 313188 25644 313240 25696
rect 445760 25644 445812 25696
rect 128268 24216 128320 24268
rect 280804 24216 280856 24268
rect 260564 24148 260616 24200
rect 431960 24148 432012 24200
rect 88248 24080 88300 24132
rect 121460 24080 121512 24132
rect 263508 24080 263560 24132
rect 500960 24080 501012 24132
rect 234436 22924 234488 22976
rect 308404 22924 308456 22976
rect 302148 22720 302200 22772
rect 442264 22720 442316 22772
rect 110328 21428 110380 21480
rect 126980 21428 127032 21480
rect 147588 21428 147640 21480
rect 169024 21428 169076 21480
rect 242716 21428 242768 21480
rect 419724 21428 419776 21480
rect 53656 21360 53708 21412
rect 111800 21360 111852 21412
rect 142068 21360 142120 21412
rect 254584 21360 254636 21412
rect 267004 21360 267056 21412
rect 498292 21360 498344 21412
rect 521016 20544 521068 20596
rect 580172 20544 580224 20596
rect 253848 19932 253900 19984
rect 462504 19932 462556 19984
rect 160008 18708 160060 18760
rect 289912 18708 289964 18760
rect 81348 18640 81400 18692
rect 118792 18640 118844 18692
rect 140688 18640 140740 18692
rect 169852 18640 169904 18692
rect 237288 18640 237340 18692
rect 401600 18640 401652 18692
rect 45376 18572 45428 18624
rect 79324 18572 79376 18624
rect 82728 18572 82780 18624
rect 147772 18572 147824 18624
rect 188896 18572 188948 18624
rect 213920 18572 213972 18624
rect 260656 18572 260708 18624
rect 494060 18572 494112 18624
rect 74448 17280 74500 17332
rect 117320 17280 117372 17332
rect 144736 17280 144788 17332
rect 169760 17280 169812 17332
rect 209688 17280 209740 17332
rect 292764 17280 292816 17332
rect 352656 17280 352708 17332
rect 396080 17280 396132 17332
rect 17868 17212 17920 17264
rect 73160 17212 73212 17264
rect 78588 17212 78640 17264
rect 146944 17212 146996 17264
rect 260748 17212 260800 17264
rect 489920 17212 489972 17264
rect 250996 15852 251048 15904
rect 455696 15852 455748 15904
rect 139308 14560 139360 14612
rect 287704 14560 287756 14612
rect 84108 14492 84160 14544
rect 89812 14492 89864 14544
rect 186964 14492 187016 14544
rect 196808 14492 196860 14544
rect 234528 14492 234580 14544
rect 390560 14492 390612 14544
rect 41328 14424 41380 14476
rect 78680 14424 78732 14476
rect 85488 14424 85540 14476
rect 119344 14424 119396 14476
rect 119896 14424 119948 14476
rect 129740 14424 129792 14476
rect 136548 14424 136600 14476
rect 168380 14424 168432 14476
rect 195244 14424 195296 14476
rect 218060 14424 218112 14476
rect 258724 14424 258776 14476
rect 480352 14424 480404 14476
rect 398104 13404 398156 13456
rect 400128 13404 400180 13456
rect 240784 13132 240836 13184
rect 409604 13132 409656 13184
rect 206928 12384 206980 12436
rect 418160 12384 418212 12436
rect 202604 12316 202656 12368
rect 416872 12316 416924 12368
rect 199844 12248 199896 12300
rect 416780 12248 416832 12300
rect 195612 12180 195664 12232
rect 415400 12180 415452 12232
rect 193036 12112 193088 12164
rect 414112 12112 414164 12164
rect 188528 12044 188580 12096
rect 414020 12044 414072 12096
rect 186136 11840 186188 11892
rect 412640 11840 412692 11892
rect 73068 11772 73120 11824
rect 87052 11772 87104 11824
rect 106188 11772 106240 11824
rect 125600 11772 125652 11824
rect 135444 11772 135496 11824
rect 400220 11772 400272 11824
rect 60648 11704 60700 11756
rect 112444 11704 112496 11756
rect 131764 11704 131816 11756
rect 398932 11704 398984 11756
rect 489920 11704 489972 11756
rect 491116 11704 491168 11756
rect 91008 11636 91060 11688
rect 92480 11636 92532 11688
rect 211068 11636 211120 11688
rect 419540 11636 419592 11688
rect 213828 11568 213880 11620
rect 419632 11568 419684 11620
rect 217968 11500 218020 11552
rect 420920 11500 420972 11552
rect 220452 11296 220504 11348
rect 422392 11296 422444 11348
rect 224776 11228 224828 11280
rect 422300 11228 422352 11280
rect 227444 11160 227496 11212
rect 423680 11160 423732 11212
rect 238668 11092 238720 11144
rect 292304 11092 292356 11144
rect 270040 11024 270092 11076
rect 282644 11024 282696 11076
rect 181996 10956 182048 11008
rect 292580 11024 292632 11076
rect 292948 11092 293000 11144
rect 426440 11092 426492 11144
rect 302516 11024 302568 11076
rect 434720 11024 434772 11076
rect 411352 10956 411404 11008
rect 177856 10752 177908 10804
rect 175188 10684 175240 10736
rect 302332 10752 302384 10804
rect 411260 10752 411312 10804
rect 170772 10616 170824 10668
rect 168288 10548 168340 10600
rect 163688 10480 163740 10532
rect 128176 10412 128228 10464
rect 292396 10480 292448 10532
rect 302332 10480 302384 10532
rect 311808 10684 311860 10736
rect 409880 10684 409932 10736
rect 408500 10616 408552 10668
rect 408592 10548 408644 10600
rect 282828 10412 282880 10464
rect 311532 10412 311584 10464
rect 407120 10480 407172 10532
rect 398840 10412 398892 10464
rect 252376 10208 252428 10260
rect 311440 10208 311492 10260
rect 311808 10208 311860 10260
rect 320180 10208 320232 10260
rect 372528 10208 372580 10260
rect 477592 10208 477644 10260
rect 255228 10140 255280 10192
rect 311624 10140 311676 10192
rect 311716 10140 311768 10192
rect 321652 10140 321704 10192
rect 372436 10140 372488 10192
rect 474556 10140 474608 10192
rect 259368 10072 259420 10124
rect 316132 10072 316184 10124
rect 369676 10072 369728 10124
rect 467472 10072 467524 10124
rect 261760 10004 261812 10056
rect 266084 9936 266136 9988
rect 317420 10004 317472 10056
rect 316040 9936 316092 9988
rect 268844 9868 268896 9920
rect 318800 9868 318852 9920
rect 273076 9664 273128 9716
rect 318892 9664 318944 9716
rect 190828 9596 190880 9648
rect 298100 9596 298152 9648
rect 314660 9596 314712 9648
rect 361488 9596 361540 9648
rect 432052 9596 432104 9648
rect 187332 9528 187384 9580
rect 296720 9528 296772 9580
rect 362868 9528 362920 9580
rect 435548 9528 435600 9580
rect 183744 9460 183796 9512
rect 180248 9392 180300 9444
rect 292396 9460 292448 9512
rect 293960 9460 294012 9512
rect 362776 9460 362828 9512
rect 439136 9460 439188 9512
rect 176660 9324 176712 9376
rect 294052 9392 294104 9444
rect 364248 9392 364300 9444
rect 442632 9392 442684 9444
rect 292672 9324 292724 9376
rect 292948 9324 293000 9376
rect 295340 9324 295392 9376
rect 365536 9324 365588 9376
rect 446220 9324 446272 9376
rect 173164 9120 173216 9172
rect 296996 9120 297048 9172
rect 366916 9120 366968 9172
rect 169576 9052 169628 9104
rect 66720 8984 66772 9036
rect 115204 8984 115256 9036
rect 166080 8984 166132 9036
rect 292856 9052 292908 9104
rect 365628 9052 365680 9104
rect 369676 9052 369728 9104
rect 369768 9052 369820 9104
rect 373724 9052 373776 9104
rect 373908 9120 373960 9172
rect 449808 9120 449860 9172
rect 456892 9052 456944 9104
rect 321560 8984 321612 9036
rect 368388 8984 368440 9036
rect 460388 8984 460440 9036
rect 21824 8916 21876 8968
rect 74540 8916 74592 8968
rect 79692 8916 79744 8968
rect 89720 8916 89772 8968
rect 102232 8916 102284 8968
rect 124312 8916 124364 8968
rect 130568 8916 130620 8968
rect 273260 8916 273312 8968
rect 273352 8916 273404 8968
rect 305092 8916 305144 8968
rect 354496 8916 354548 8968
rect 393320 8916 393372 8968
rect 393412 8916 393464 8968
rect 463976 8916 464028 8968
rect 194416 8848 194468 8900
rect 299572 8848 299624 8900
rect 360108 8848 360160 8900
rect 428464 8848 428516 8900
rect 197912 8780 197964 8832
rect 299480 8780 299532 8832
rect 360016 8780 360068 8832
rect 424968 8780 425020 8832
rect 201500 8576 201552 8628
rect 300860 8576 300912 8628
rect 358728 8576 358780 8628
rect 421380 8576 421432 8628
rect 205088 8508 205140 8560
rect 302240 8508 302292 8560
rect 357348 8508 357400 8560
rect 417884 8508 417936 8560
rect 208584 8440 208636 8492
rect 302424 8440 302476 8492
rect 357256 8440 357308 8492
rect 414296 8440 414348 8492
rect 212172 8372 212224 8424
rect 303620 8372 303672 8424
rect 355968 8372 356020 8424
rect 410800 8372 410852 8424
rect 215668 8304 215720 8356
rect 305000 8304 305052 8356
rect 354588 8304 354640 8356
rect 407212 8304 407264 8356
rect 219256 8236 219308 8288
rect 248880 8236 248932 8288
rect 430856 8236 430908 8288
rect 245568 8032 245620 8084
rect 434444 8032 434496 8084
rect 246948 7964 247000 8016
rect 437940 7964 437992 8016
rect 248328 7896 248380 7948
rect 441528 7896 441580 7948
rect 248236 7828 248288 7880
rect 445024 7828 445076 7880
rect 251088 7760 251140 7812
rect 245476 7692 245528 7744
rect 448612 7760 448664 7812
rect 452108 7692 452160 7744
rect 244188 7488 244240 7540
rect 427268 7488 427320 7540
rect 242808 7420 242860 7472
rect 412640 7420 412692 7472
rect 412732 7420 412784 7472
rect 577412 7420 577464 7472
rect 249708 7352 249760 7404
rect 284208 7352 284260 7404
rect 367008 7352 367060 7404
rect 453304 7352 453356 7404
rect 471060 7352 471112 7404
rect 394516 7284 394568 7336
rect 398656 7284 398708 7336
rect 398748 7284 398800 7336
rect 397368 7216 397420 7268
rect 573916 7284 573968 7336
rect 397276 7148 397328 7200
rect 570328 7216 570380 7268
rect 408316 7148 408368 7200
rect 408408 7148 408460 7200
rect 566832 7148 566884 7200
rect 395988 6944 396040 6996
rect 398840 6944 398892 6996
rect 398932 6944 398984 6996
rect 563244 6944 563296 6996
rect 371148 6876 371200 6928
rect 293684 6808 293736 6860
rect 324412 6808 324464 6860
rect 290188 6740 290240 6792
rect 324320 6740 324372 6792
rect 325608 6740 325660 6792
rect 332600 6740 332652 6792
rect 286600 6672 286652 6724
rect 322940 6672 322992 6724
rect 323032 6672 323084 6724
rect 331312 6672 331364 6724
rect 223488 6604 223540 6656
rect 345756 6808 345808 6860
rect 346216 6808 346268 6860
rect 375288 6808 375340 6860
rect 386236 6808 386288 6860
rect 531320 6808 531372 6860
rect 347688 6740 347740 6792
rect 378876 6740 378928 6792
rect 388996 6740 389048 6792
rect 534908 6740 534960 6792
rect 340788 6672 340840 6724
rect 348976 6672 349028 6724
rect 382372 6672 382424 6724
rect 389088 6672 389140 6724
rect 538404 6672 538456 6724
rect 340696 6604 340748 6656
rect 348792 6604 348844 6656
rect 349068 6604 349120 6656
rect 385960 6604 386012 6656
rect 390468 6604 390520 6656
rect 394608 6604 394660 6656
rect 541992 6604 542044 6656
rect 223396 6400 223448 6452
rect 349252 6400 349304 6452
rect 350356 6400 350408 6452
rect 350448 6400 350500 6452
rect 389456 6400 389508 6452
rect 391756 6400 391808 6452
rect 545488 6400 545540 6452
rect 224868 6332 224920 6384
rect 184848 6264 184900 6316
rect 193220 6264 193272 6316
rect 226156 6264 226208 6316
rect 351828 6332 351880 6384
rect 352840 6264 352892 6316
rect 387708 6264 387760 6316
rect 391848 6332 391900 6384
rect 549076 6332 549128 6384
rect 76196 6196 76248 6248
rect 88340 6196 88392 6248
rect 98644 6196 98696 6248
rect 124220 6196 124272 6248
rect 188988 6196 189040 6248
rect 210976 6196 211028 6248
rect 226248 6196 226300 6248
rect 359924 6196 359976 6248
rect 380808 6196 380860 6248
rect 393044 6264 393096 6316
rect 393228 6264 393280 6316
rect 394608 6196 394660 6248
rect 552664 6264 552716 6316
rect 463884 6239 463936 6248
rect 463884 6205 463893 6239
rect 463893 6205 463927 6239
rect 463927 6205 463936 6239
rect 463884 6196 463936 6205
rect 556160 6196 556212 6248
rect 26516 6128 26568 6180
rect 75920 6128 75972 6180
rect 77392 6128 77444 6180
rect 118700 6128 118752 6180
rect 125876 6128 125928 6180
rect 165620 6128 165672 6180
rect 191656 6128 191708 6180
rect 221556 6128 221608 6180
rect 227628 6128 227680 6180
rect 363512 6128 363564 6180
rect 379428 6128 379480 6180
rect 502156 6128 502208 6180
rect 559748 6128 559800 6180
rect 297272 6060 297324 6112
rect 325700 6060 325752 6112
rect 346308 6060 346360 6112
rect 371700 6060 371752 6112
rect 386144 6060 386196 6112
rect 527824 6060 527876 6112
rect 300768 5856 300820 5908
rect 327080 5856 327132 5908
rect 344928 5856 344980 5908
rect 368204 5856 368256 5908
rect 384948 5856 385000 5908
rect 524236 5856 524288 5908
rect 304356 5788 304408 5840
rect 327172 5788 327224 5840
rect 331220 5788 331272 5840
rect 337936 5788 337988 5840
rect 343364 5788 343416 5840
rect 343548 5788 343600 5840
rect 364616 5788 364668 5840
rect 383568 5788 383620 5840
rect 520740 5788 520792 5840
rect 520924 5788 520976 5840
rect 580172 5788 580224 5840
rect 307944 5720 307996 5772
rect 328460 5720 328512 5772
rect 339408 5720 339460 5772
rect 315028 5652 315080 5704
rect 282828 5584 282880 5636
rect 311440 5584 311492 5636
rect 329840 5652 329892 5704
rect 343456 5720 343508 5772
rect 361120 5720 361172 5772
rect 383476 5720 383528 5772
rect 517152 5720 517204 5772
rect 346952 5652 347004 5704
rect 86868 5516 86920 5568
rect 91100 5516 91152 5568
rect 184204 5516 184256 5568
rect 189724 5516 189776 5568
rect 275928 5516 275980 5568
rect 316040 5516 316092 5568
rect 318524 5516 318576 5568
rect 329196 5584 329248 5636
rect 334072 5584 334124 5636
rect 334164 5584 334216 5636
rect 329932 5516 329984 5568
rect 332692 5516 332744 5568
rect 333980 5516 334032 5568
rect 338028 5584 338080 5636
rect 339868 5584 339920 5636
rect 342168 5584 342220 5636
rect 357532 5652 357584 5704
rect 382188 5652 382240 5704
rect 513564 5652 513616 5704
rect 356336 5584 356388 5636
rect 380716 5584 380768 5636
rect 510068 5584 510120 5636
rect 383660 5516 383712 5568
rect 499672 5516 499724 5568
rect 499764 5516 499816 5568
rect 514576 5516 514628 5568
rect 63224 5312 63276 5364
rect 114560 5312 114612 5364
rect 200028 5312 200080 5364
rect 257068 5312 257120 5364
rect 274456 5312 274508 5364
rect 277124 5312 277176 5364
rect 56048 5244 56100 5296
rect 113272 5244 113324 5296
rect 201408 5244 201460 5296
rect 205272 5244 205324 5296
rect 205548 5244 205600 5296
rect 267740 5244 267792 5296
rect 274548 5244 274600 5296
rect 48964 5176 49016 5228
rect 110420 5176 110472 5228
rect 202788 5176 202840 5228
rect 205364 5176 205416 5228
rect 205456 5176 205508 5228
rect 271236 5176 271288 5228
rect 271788 5176 271840 5228
rect 278688 5312 278740 5364
rect 544384 5312 544436 5364
rect 282828 5244 282880 5296
rect 547880 5244 547932 5296
rect 1676 5108 1728 5160
rect 70400 5108 70452 5160
rect 97908 5108 97960 5160
rect 108120 5108 108172 5160
rect 191748 5108 191800 5160
rect 219440 5108 219492 5160
rect 274824 5108 274876 5160
rect 277216 5108 277268 5160
rect 551468 5176 551520 5228
rect 2872 5040 2924 5092
rect 71780 5040 71832 5092
rect 99196 5040 99248 5092
rect 115204 5040 115256 5092
rect 193128 5040 193180 5092
rect 278320 5040 278372 5092
rect 554964 5108 555016 5160
rect 558552 5040 558604 5092
rect 572 4972 624 5024
rect 70492 4972 70544 5024
rect 100668 4972 100720 5024
rect 118792 4972 118844 5024
rect 204168 4972 204220 5024
rect 209688 4972 209740 5024
rect 260656 4972 260708 5024
rect 266268 4972 266320 5024
rect 509240 4972 509292 5024
rect 562048 4972 562100 5024
rect 4068 4768 4120 4820
rect 100760 4768 100812 4820
rect 102048 4768 102100 4820
rect 122288 4768 122340 4820
rect 202696 4768 202748 4820
rect 209596 4768 209648 4820
rect 264152 4768 264204 4820
rect 266176 4768 266228 4820
rect 480260 4768 480312 4820
rect 480352 4768 480404 4820
rect 489828 4768 489880 4820
rect 489920 4768 489972 4820
rect 499396 4768 499448 4820
rect 499488 4768 499540 4820
rect 565636 4768 565688 4820
rect 47860 4700 47912 4752
rect 81440 4700 81492 4752
rect 99288 4700 99340 4752
rect 111616 4700 111668 4752
rect 199936 4700 199988 4752
rect 253480 4700 253532 4752
rect 271696 4700 271748 4752
rect 51356 4632 51408 4684
rect 81532 4632 81584 4684
rect 96160 4632 96212 4684
rect 104532 4632 104584 4684
rect 198648 4632 198700 4684
rect 249984 4632 250036 4684
rect 54944 4564 54996 4616
rect 82820 4564 82872 4616
rect 197268 4564 197320 4616
rect 246396 4564 246448 4616
rect 273168 4564 273220 4616
rect 540796 4700 540848 4752
rect 537208 4632 537260 4684
rect 533712 4564 533764 4616
rect 65524 4496 65576 4548
rect 85580 4496 85632 4548
rect 197176 4496 197228 4548
rect 242900 4496 242952 4548
rect 270408 4496 270460 4548
rect 530124 4496 530176 4548
rect 69112 4428 69164 4480
rect 86960 4428 87012 4480
rect 195888 4428 195940 4480
rect 239312 4428 239364 4480
rect 268936 4428 268988 4480
rect 526628 4428 526680 4480
rect 96436 4224 96488 4276
rect 101036 4224 101088 4276
rect 194232 4224 194284 4276
rect 235724 4224 235776 4276
rect 269028 4224 269080 4276
rect 523040 4224 523092 4276
rect 95148 4156 95200 4208
rect 97448 4156 97500 4208
rect 135352 4156 135404 4208
rect 194324 4156 194376 4208
rect 232228 4156 232280 4208
rect 267648 4156 267700 4208
rect 519544 4156 519596 4208
rect 6460 4088 6512 4140
rect 7564 4088 7616 4140
rect 85672 4088 85724 4140
rect 149060 4088 149112 4140
rect 158904 4088 158956 4140
rect 160008 4088 160060 4140
rect 164884 4088 164936 4140
rect 165528 4088 165580 4140
rect 228732 4088 228784 4140
rect 273628 4088 273680 4140
rect 274364 4088 274416 4140
rect 277216 4088 277268 4140
rect 278044 4088 278096 4140
rect 283104 4088 283156 4140
rect 284208 4088 284260 4140
rect 284300 4088 284352 4140
rect 285588 4088 285640 4140
rect 287796 4088 287848 4140
rect 288348 4088 288400 4140
rect 291384 4088 291436 4140
rect 292488 4088 292540 4140
rect 298468 4088 298520 4140
rect 299388 4088 299440 4140
rect 305552 4088 305604 4140
rect 308496 4088 308548 4140
rect 309048 4088 309100 4140
rect 309784 4088 309836 4140
rect 14740 4020 14792 4072
rect 18604 4020 18656 4072
rect 46664 4020 46716 4072
rect 132960 4020 133012 4072
rect 133788 4020 133840 4072
rect 134156 4020 134208 4072
rect 135168 4020 135220 4072
rect 280068 4020 280120 4072
rect 383660 4088 383712 4140
rect 387156 4088 387208 4140
rect 461216 4088 461268 4140
rect 468024 4088 468076 4140
rect 383568 4020 383620 4072
rect 461124 4020 461176 4072
rect 462412 4020 462464 4072
rect 469220 4020 469272 4072
rect 470692 4020 470744 4072
rect 510528 4088 510580 4140
rect 553768 4088 553820 4140
rect 509148 4020 509200 4072
rect 557356 4020 557408 4072
rect 43076 3952 43128 4004
rect 138112 3952 138164 4004
rect 157800 3952 157852 4004
rect 173900 3952 173952 4004
rect 333888 3952 333940 4004
rect 336004 3952 336056 4004
rect 379980 3952 380032 4004
rect 460572 3952 460624 4004
rect 460848 3952 460900 4004
rect 483204 3952 483256 4004
rect 489184 3952 489236 4004
rect 492312 3952 492364 4004
rect 498016 3952 498068 4004
rect 515956 3952 516008 4004
rect 560852 3952 560904 4004
rect 39580 3884 39632 3936
rect 138020 3884 138072 3936
rect 154212 3884 154264 3936
rect 172612 3884 172664 3936
rect 186044 3884 186096 3936
rect 203892 3884 203944 3936
rect 276020 3884 276072 3936
rect 277308 3884 277360 3936
rect 376484 3884 376536 3936
rect 451372 3884 451424 3936
rect 455512 3884 455564 3936
rect 460664 3884 460716 3936
rect 480628 3884 480680 3936
rect 496728 3884 496780 3936
rect 507676 3884 507728 3936
rect 509056 3884 509108 3936
rect 564440 3884 564492 3936
rect 35992 3680 36044 3732
rect 116400 3680 116452 3732
rect 117228 3680 117280 3732
rect 117596 3680 117648 3732
rect 124680 3680 124732 3732
rect 158720 3680 158772 3732
rect 168380 3680 168432 3732
rect 176016 3680 176068 3732
rect 187608 3680 187660 3732
rect 207388 3680 207440 3732
rect 226340 3680 226392 3732
rect 227536 3680 227588 3732
rect 251180 3680 251232 3732
rect 252376 3680 252428 3732
rect 319720 3680 319772 3732
rect 320824 3680 320876 3732
rect 358728 3680 358780 3732
rect 451280 3680 451332 3732
rect 454408 3680 454460 3732
rect 454500 3680 454552 3732
rect 455328 3680 455380 3732
rect 477684 3680 477736 3732
rect 495348 3680 495400 3732
rect 500592 3680 500644 3732
rect 32496 3612 32548 3664
rect 8760 3544 8812 3596
rect 14464 3544 14516 3596
rect 15936 3544 15988 3596
rect 19984 3544 20036 3596
rect 27712 3544 27764 3596
rect 28908 3544 28960 3596
rect 31300 3544 31352 3596
rect 32404 3544 32456 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 136640 3612 136692 3664
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 7656 3408 7708 3460
rect 10324 3408 10376 3460
rect 19432 3408 19484 3460
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 126980 3476 127032 3528
rect 128268 3476 128320 3528
rect 133972 3544 134024 3596
rect 134064 3544 134116 3596
rect 158812 3612 158864 3664
rect 160100 3612 160152 3664
rect 405740 3612 405792 3664
rect 415492 3612 415544 3664
rect 416688 3612 416740 3664
rect 422576 3612 422628 3664
rect 423588 3612 423640 3664
rect 473544 3612 473596 3664
rect 498108 3612 498160 3664
rect 511264 3680 511316 3732
rect 511816 3680 511868 3732
rect 516232 3680 516284 3732
rect 514760 3612 514812 3664
rect 516048 3612 516100 3664
rect 518624 3680 518676 3732
rect 568028 3680 568080 3732
rect 139400 3544 139452 3596
rect 143540 3544 143592 3596
rect 144736 3544 144788 3596
rect 156604 3544 156656 3596
rect 405832 3544 405884 3596
rect 411904 3544 411956 3596
rect 470784 3544 470836 3596
rect 485044 3544 485096 3596
rect 489920 3544 489972 3596
rect 491208 3544 491260 3596
rect 499304 3544 499356 3596
rect 518348 3544 518400 3596
rect 571524 3612 571576 3664
rect 138848 3476 138900 3528
rect 139308 3476 139360 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 150624 3476 150676 3528
rect 151728 3476 151780 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 155408 3476 155460 3528
rect 155868 3476 155920 3528
rect 404360 3476 404412 3528
rect 408408 3476 408460 3528
rect 470600 3476 470652 3528
rect 479340 3476 479392 3528
rect 480168 3476 480220 3528
rect 135260 3408 135312 3460
rect 149520 3408 149572 3460
rect 402980 3408 403032 3460
rect 404820 3408 404872 3460
rect 461584 3408 461636 3460
rect 462228 3408 462280 3460
rect 462320 3408 462372 3460
rect 467932 3408 467984 3460
rect 468668 3408 468720 3460
rect 469128 3408 469180 3460
rect 486424 3476 486476 3528
rect 487068 3476 487120 3528
rect 487804 3476 487856 3528
rect 493968 3476 494020 3528
rect 497096 3476 497148 3528
rect 500776 3476 500828 3528
rect 521844 3476 521896 3528
rect 575112 3544 575164 3596
rect 579804 3476 579856 3528
rect 28908 3340 28960 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 41880 3340 41932 3392
rect 42708 3340 42760 3392
rect 44272 3340 44324 3392
rect 45376 3340 45428 3392
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 52552 3340 52604 3392
rect 53656 3340 53708 3392
rect 57244 3340 57296 3392
rect 57888 3340 57940 3392
rect 58440 3340 58492 3392
rect 59268 3340 59320 3392
rect 59636 3340 59688 3392
rect 60648 3340 60700 3392
rect 60832 3340 60884 3392
rect 61936 3340 61988 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 67916 3340 67968 3392
rect 68928 3340 68980 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 75000 3340 75052 3392
rect 75828 3340 75880 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 82084 3340 82136 3392
rect 82728 3340 82780 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 84476 3340 84528 3392
rect 85488 3340 85540 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 91560 3340 91612 3392
rect 92388 3340 92440 3392
rect 150532 3340 150584 3392
rect 153016 3340 153068 3392
rect 167184 3340 167236 3392
rect 168288 3340 168340 3392
rect 174268 3340 174320 3392
rect 175188 3340 175240 3392
rect 175464 3340 175516 3392
rect 178132 3340 178184 3392
rect 181444 3340 181496 3392
rect 181996 3340 182048 3392
rect 184940 3340 184992 3392
rect 186136 3340 186188 3392
rect 206192 3340 206244 3392
rect 206928 3340 206980 3392
rect 209780 3340 209832 3392
rect 211068 3340 211120 3392
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 216864 3340 216916 3392
rect 217968 3340 218020 3392
rect 222752 3340 222804 3392
rect 223304 3340 223356 3392
rect 223948 3340 224000 3392
rect 224776 3340 224828 3392
rect 229836 3340 229888 3392
rect 230388 3340 230440 3392
rect 231032 3340 231084 3392
rect 231676 3340 231728 3392
rect 233424 3340 233476 3392
rect 234436 3340 234488 3392
rect 234620 3340 234672 3392
rect 235816 3340 235868 3392
rect 238116 3340 238168 3392
rect 238668 3340 238720 3392
rect 240508 3340 240560 3392
rect 241428 3340 241480 3392
rect 241704 3340 241756 3392
rect 242624 3340 242676 3392
rect 247592 3340 247644 3392
rect 248144 3340 248196 3392
rect 248788 3340 248840 3392
rect 249616 3340 249668 3392
rect 254676 3340 254728 3392
rect 255228 3340 255280 3392
rect 255872 3340 255924 3392
rect 256424 3340 256476 3392
rect 259460 3340 259512 3392
rect 260564 3340 260616 3392
rect 265348 3340 265400 3392
rect 266084 3340 266136 3392
rect 266544 3340 266596 3392
rect 267556 3340 267608 3392
rect 272432 3340 272484 3392
rect 273076 3340 273128 3392
rect 312636 3340 312688 3392
rect 313188 3340 313240 3392
rect 316224 3340 316276 3392
rect 318064 3340 318116 3392
rect 323308 3340 323360 3392
rect 324228 3340 324280 3392
rect 330392 3340 330444 3392
rect 331128 3340 331180 3392
rect 335360 3340 335412 3392
rect 336280 3340 336332 3392
rect 337476 3340 337528 3392
rect 338764 3340 338816 3392
rect 348056 3340 348108 3392
rect 349804 3340 349856 3392
rect 351644 3340 351696 3392
rect 352564 3340 352616 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 390652 3340 390704 3392
rect 463700 3340 463752 3392
rect 495900 3408 495952 3460
rect 500868 3408 500920 3460
rect 518992 3408 519044 3460
rect 583392 3408 583444 3460
rect 499396 3340 499448 3392
rect 507768 3340 507820 3392
rect 550272 3340 550324 3392
rect 89168 3136 89220 3188
rect 92756 3136 92808 3188
rect 150440 3136 150492 3188
rect 171968 3136 172020 3188
rect 175924 3136 175976 3188
rect 182088 3136 182140 3188
rect 186136 3136 186188 3188
rect 199108 3136 199160 3188
rect 199844 3136 199896 3188
rect 322112 3136 322164 3188
rect 322848 3136 322900 3188
rect 390560 3136 390612 3188
rect 391848 3136 391900 3188
rect 394240 3136 394292 3188
rect 17040 3068 17092 3120
rect 17868 3068 17920 3120
rect 99840 3068 99892 3120
rect 153200 3068 153252 3120
rect 397736 3068 397788 3120
rect 460848 3068 460900 3120
rect 13544 3000 13596 3052
rect 15844 3000 15896 3052
rect 103336 3000 103388 3052
rect 153292 3000 153344 3052
rect 340972 3000 341024 3052
rect 344284 3000 344336 3052
rect 355232 3000 355284 3052
rect 358084 3000 358136 3052
rect 401324 3000 401376 3052
rect 461308 3136 461360 3188
rect 465080 3136 465132 3188
rect 465172 3136 465224 3188
rect 466368 3136 466420 3188
rect 472256 3136 472308 3188
rect 473268 3136 473320 3188
rect 506388 3136 506440 3188
rect 546684 3136 546736 3188
rect 465356 3068 465408 3120
rect 506296 3068 506348 3120
rect 543188 3068 543240 3120
rect 466460 3000 466512 3052
rect 505008 3000 505060 3052
rect 539600 3000 539652 3052
rect 105728 2932 105780 2984
rect 106188 2932 106240 2984
rect 106924 2932 106976 2984
rect 107568 2932 107620 2984
rect 109316 2932 109368 2984
rect 110328 2932 110380 2984
rect 110512 2932 110564 2984
rect 155960 2932 156012 2984
rect 192024 2932 192076 2984
rect 193036 2932 193088 2984
rect 258264 2932 258316 2984
rect 259368 2932 259420 2984
rect 415492 2932 415544 2984
rect 416596 2932 416648 2984
rect 418988 2932 419040 2984
rect 426164 2932 426216 2984
rect 474832 2932 474884 2984
rect 503628 2932 503680 2984
rect 536104 2932 536156 2984
rect 73804 2864 73856 2916
rect 74448 2864 74500 2916
rect 114008 2864 114060 2916
rect 156052 2864 156104 2916
rect 280712 2864 280764 2916
rect 281448 2864 281500 2916
rect 429660 2864 429712 2916
rect 476120 2864 476172 2916
rect 503536 2864 503588 2916
rect 532516 2864 532568 2916
rect 128360 2796 128412 2848
rect 132224 2796 132276 2848
rect 157340 2796 157392 2848
rect 433248 2796 433300 2848
rect 436744 2796 436796 2848
rect 437388 2796 437440 2848
rect 476212 2796 476264 2848
rect 502064 2796 502116 2848
rect 529020 2796 529072 2848
rect 440332 2592 440384 2644
rect 441712 2592 441764 2644
rect 447416 2592 447468 2644
rect 525432 2592 525484 2644
rect 121092 2524 121144 2576
rect 340880 1980 340932 2032
rect 342168 1980 342220 2032
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 680338 3464 697303
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 680332 3476 680338
rect 3424 680274 3476 680280
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 658170 3464 671191
rect 3528 669322 3556 684247
rect 8220 682446 8248 702406
rect 24320 699718 24348 703520
rect 40512 700534 40540 703520
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 41328 700528 41380 700534
rect 41328 700470 41380 700476
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 682514 24808 699654
rect 41340 682582 41368 700470
rect 56796 700330 56824 703520
rect 72988 702434 73016 703520
rect 72988 702406 73108 702434
rect 56784 700324 56836 700330
rect 56784 700266 56836 700272
rect 57888 700324 57940 700330
rect 57888 700266 57940 700272
rect 57900 682650 57928 700266
rect 57888 682644 57940 682650
rect 57888 682586 57940 682592
rect 41328 682576 41380 682582
rect 41328 682518 41380 682524
rect 24768 682508 24820 682514
rect 24768 682450 24820 682456
rect 73080 682446 73108 702406
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 121656 699718 121684 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154528 702434
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 89640 682514 89668 699654
rect 106200 682582 106228 699654
rect 108396 682644 108448 682650
rect 108396 682586 108448 682592
rect 95608 682576 95660 682582
rect 95608 682518 95660 682524
rect 106188 682576 106240 682582
rect 106188 682518 106240 682524
rect 82820 682508 82872 682514
rect 82820 682450 82872 682456
rect 89628 682508 89680 682514
rect 89628 682450 89680 682456
rect 8208 682440 8260 682446
rect 8208 682382 8260 682388
rect 71044 682440 71096 682446
rect 71044 682382 71096 682388
rect 73068 682440 73120 682446
rect 73068 682382 73120 682388
rect 66996 680332 67048 680338
rect 66996 680274 67048 680280
rect 67008 679153 67036 680274
rect 71056 680218 71084 682382
rect 82832 680218 82860 682450
rect 95620 680218 95648 682518
rect 108408 680218 108436 682586
rect 122760 682446 122788 699654
rect 137940 682514 137968 702406
rect 154500 682582 154528 702406
rect 170324 699718 170352 703520
rect 186516 700330 186544 703520
rect 186504 700324 186556 700330
rect 186504 700266 186556 700272
rect 187608 700324 187660 700330
rect 187608 700266 187660 700272
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 146852 682576 146904 682582
rect 146852 682518 146904 682524
rect 154488 682576 154540 682582
rect 154488 682518 154540 682524
rect 134064 682508 134116 682514
rect 134064 682450 134116 682456
rect 137928 682508 137980 682514
rect 137928 682450 137980 682456
rect 121184 682440 121236 682446
rect 121184 682382 121236 682388
rect 122748 682440 122800 682446
rect 122748 682382 122800 682388
rect 121196 680218 121224 682382
rect 134076 680218 134104 682450
rect 146864 680218 146892 682518
rect 171060 682446 171088 699654
rect 185216 682576 185268 682582
rect 185216 682518 185268 682524
rect 172428 682508 172480 682514
rect 172428 682450 172480 682456
rect 159640 682440 159692 682446
rect 159640 682382 159692 682388
rect 171048 682440 171100 682446
rect 171048 682382 171100 682388
rect 159652 680218 159680 682382
rect 172440 680218 172468 682450
rect 185228 680218 185256 682518
rect 187620 682514 187648 700266
rect 187608 682508 187660 682514
rect 187608 682450 187660 682456
rect 202800 682446 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 219360 682514 219388 702406
rect 235184 699718 235212 703520
rect 251468 699718 251496 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 251456 699712 251508 699718
rect 251456 699654 251508 699660
rect 252468 699712 252520 699718
rect 252468 699654 252520 699660
rect 210792 682508 210844 682514
rect 210792 682450 210844 682456
rect 219348 682508 219400 682514
rect 219348 682450 219400 682456
rect 198004 682440 198056 682446
rect 198004 682382 198056 682388
rect 202788 682440 202840 682446
rect 202788 682382 202840 682388
rect 198016 680218 198044 682382
rect 210804 680218 210832 682450
rect 235920 682446 235948 699654
rect 236368 682508 236420 682514
rect 236368 682450 236420 682456
rect 223580 682440 223632 682446
rect 223580 682382 223632 682388
rect 235908 682440 235960 682446
rect 235908 682382 235960 682388
rect 223592 680218 223620 682382
rect 236380 680218 236408 682450
rect 252480 682446 252508 699654
rect 267660 682446 267688 703520
rect 283852 702434 283880 703520
rect 283852 702406 284248 702434
rect 284220 682922 284248 702406
rect 300136 699718 300164 703520
rect 316328 699718 316356 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 364996 700330 365024 703520
rect 378048 700392 378100 700398
rect 378048 700334 378100 700340
rect 339408 700324 339460 700330
rect 339408 700266 339460 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 351828 700324 351880 700330
rect 351828 700266 351880 700272
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 365628 700324 365680 700330
rect 365628 700266 365680 700272
rect 299480 699712 299532 699718
rect 299480 699654 299532 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 313188 699712 313240 699718
rect 313188 699654 313240 699660
rect 316316 699712 316368 699718
rect 316316 699654 316368 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 284208 682916 284260 682922
rect 284208 682858 284260 682864
rect 287612 682916 287664 682922
rect 287612 682858 287664 682864
rect 249248 682440 249300 682446
rect 249248 682382 249300 682388
rect 252468 682440 252520 682446
rect 252468 682382 252520 682388
rect 262036 682440 262088 682446
rect 262036 682382 262088 682388
rect 267648 682440 267700 682446
rect 267648 682382 267700 682388
rect 274824 682440 274876 682446
rect 274824 682382 274876 682388
rect 249260 680218 249288 682382
rect 262048 680218 262076 682382
rect 274836 680218 274864 682382
rect 287624 680218 287652 682858
rect 71044 680190 71084 680218
rect 82820 680190 82860 680218
rect 95608 680190 95648 680218
rect 108396 680190 108436 680218
rect 121184 680190 121224 680218
rect 134064 680190 134104 680218
rect 146852 680190 146892 680218
rect 159640 680190 159680 680218
rect 172428 680190 172468 680218
rect 185216 680190 185256 680218
rect 198004 680190 198044 680218
rect 210792 680190 210832 680218
rect 223580 680190 223620 680218
rect 236368 680190 236408 680218
rect 249248 680190 249288 680218
rect 262036 680190 262076 680218
rect 274824 680190 274864 680218
rect 287612 680190 287652 680218
rect 71044 680000 71072 680190
rect 82820 680000 82848 680190
rect 95608 680000 95636 680190
rect 108396 680000 108424 680190
rect 121184 680000 121212 680190
rect 134064 680000 134092 680190
rect 146852 680000 146880 680190
rect 159640 680000 159668 680190
rect 172428 680000 172456 680190
rect 185216 680000 185244 680190
rect 198004 680000 198032 680190
rect 210792 680000 210820 680190
rect 223580 680000 223608 680190
rect 236368 680000 236396 680190
rect 249248 680000 249276 680190
rect 262036 680000 262064 680190
rect 274824 680000 274852 680190
rect 287612 680000 287640 680190
rect 299492 680082 299520 699654
rect 313200 680218 313228 699654
rect 327000 681766 327028 699654
rect 339420 681766 339448 700266
rect 325976 681760 326028 681766
rect 325976 681702 326028 681708
rect 326988 681760 327040 681766
rect 326988 681702 327040 681708
rect 338764 681760 338816 681766
rect 338764 681702 338816 681708
rect 339408 681760 339460 681766
rect 339408 681702 339460 681708
rect 325988 680218 326016 681702
rect 338776 680218 338804 681702
rect 313188 680190 313228 680218
rect 325976 680190 326016 680218
rect 338764 680190 338804 680218
rect 299492 680054 300428 680082
rect 300400 680000 300428 680054
rect 313188 680000 313216 680190
rect 325976 680000 326004 680190
rect 338764 680000 338792 680190
rect 351840 680082 351868 700266
rect 365640 681766 365668 700266
rect 378060 681766 378088 700334
rect 381188 700330 381216 703520
rect 397472 700398 397500 703520
rect 402888 700460 402940 700466
rect 402888 700402 402940 700408
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 381176 700324 381228 700330
rect 381176 700266 381228 700272
rect 390468 700324 390520 700330
rect 390468 700266 390520 700272
rect 390480 681766 390508 700266
rect 364432 681760 364484 681766
rect 364432 681702 364484 681708
rect 365628 681760 365680 681766
rect 365628 681702 365680 681708
rect 377220 681760 377272 681766
rect 377220 681702 377272 681708
rect 378048 681760 378100 681766
rect 378048 681702 378100 681708
rect 390008 681760 390060 681766
rect 390008 681702 390060 681708
rect 390468 681760 390520 681766
rect 390468 681702 390520 681708
rect 364444 680218 364472 681702
rect 377232 680218 377260 681702
rect 390020 680218 390048 681702
rect 351552 680054 351868 680082
rect 364432 680190 364472 680218
rect 377220 680190 377260 680218
rect 390008 680190 390048 680218
rect 351552 680000 351580 680054
rect 364432 680000 364460 680190
rect 377220 680000 377248 680190
rect 390008 680000 390036 680190
rect 402900 680082 402928 700402
rect 413664 700330 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 441528 700460 441580 700466
rect 441528 700402 441580 700408
rect 416688 700392 416740 700398
rect 416688 700334 416740 700340
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 416700 681766 416728 700334
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 681766 429148 700266
rect 415584 681760 415636 681766
rect 415584 681702 415636 681708
rect 416688 681760 416740 681766
rect 416688 681702 416740 681708
rect 428372 681760 428424 681766
rect 428372 681702 428424 681708
rect 429108 681760 429160 681766
rect 429108 681702 429160 681708
rect 415596 680218 415624 681702
rect 428384 680218 428412 681702
rect 402796 680054 402928 680082
rect 415584 680190 415624 680218
rect 428372 680190 428412 680218
rect 402796 680000 402824 680054
rect 415584 680000 415612 680190
rect 428372 680000 428400 680190
rect 441540 680082 441568 700402
rect 446140 700398 446168 703520
rect 446128 700392 446180 700398
rect 446128 700334 446180 700340
rect 453948 700392 454000 700398
rect 453948 700334 454000 700340
rect 453960 680218 453988 700334
rect 462332 700330 462360 703520
rect 478524 700466 478552 703520
rect 480168 700528 480220 700534
rect 480168 700470 480220 700476
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 467748 700324 467800 700330
rect 467748 700266 467800 700272
rect 467760 681766 467788 700266
rect 480180 681766 480208 700470
rect 492588 700460 492640 700466
rect 492588 700402 492640 700408
rect 466736 681760 466788 681766
rect 466736 681702 466788 681708
rect 467748 681760 467800 681766
rect 467748 681702 467800 681708
rect 479616 681760 479668 681766
rect 479616 681702 479668 681708
rect 480168 681760 480220 681766
rect 480168 681702 480220 681708
rect 466748 680218 466776 681702
rect 479628 680218 479656 681702
rect 441160 680054 441568 680082
rect 453948 680190 453988 680218
rect 466736 680190 466776 680218
rect 479616 680190 479656 680218
rect 441160 680000 441188 680054
rect 453948 680000 453976 680190
rect 466736 680000 466764 680190
rect 479616 680000 479644 680190
rect 492600 680082 492628 700402
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 506388 700392 506440 700398
rect 506388 700334 506440 700340
rect 506400 681766 506428 700334
rect 511000 700330 511028 703520
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 575860 700330 575888 703520
rect 510988 700324 511040 700330
rect 510988 700266 511040 700272
rect 517428 700324 517480 700330
rect 517428 700266 517480 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 505192 681760 505244 681766
rect 505192 681702 505244 681708
rect 506388 681760 506440 681766
rect 506388 681702 506440 681708
rect 505204 680218 505232 681702
rect 492404 680054 492628 680082
rect 505192 680190 505232 680218
rect 492404 680000 492432 680054
rect 505192 680000 505220 680190
rect 517440 680082 517468 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 520924 696992 520976 696998
rect 520924 696934 520976 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 517060 680054 517468 680082
rect 517060 680000 517088 680054
rect 66994 679144 67050 679153
rect 66994 679079 67050 679088
rect 520936 678881 520964 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 521016 683188 521068 683194
rect 521016 683130 521068 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 520922 678872 520978 678881
rect 520922 678807 520978 678816
rect 520924 670880 520976 670886
rect 520924 670822 520976 670828
rect 3516 669316 3568 669322
rect 3516 669258 3568 669264
rect 67180 669316 67232 669322
rect 67180 669258 67232 669264
rect 67192 668953 67220 669258
rect 67178 668944 67234 668953
rect 67178 668879 67234 668888
rect 3514 658200 3570 658209
rect 3424 658164 3476 658170
rect 3514 658135 3570 658144
rect 67364 658164 67416 658170
rect 3424 658106 3476 658112
rect 3528 647222 3556 658135
rect 67364 658106 67416 658112
rect 67376 657801 67404 658106
rect 67362 657792 67418 657801
rect 67362 657727 67418 657736
rect 520936 657257 520964 670822
rect 521028 668545 521056 683130
rect 580172 670880 580224 670886
rect 580172 670822 580224 670828
rect 580184 670721 580212 670822
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 521014 668536 521070 668545
rect 521014 668471 521070 668480
rect 580170 657384 580226 657393
rect 580170 657319 580226 657328
rect 520922 657248 520978 657257
rect 520922 657183 520978 657192
rect 580184 656946 580212 657319
rect 521016 656940 521068 656946
rect 521016 656882 521068 656888
rect 580172 656940 580224 656946
rect 580172 656882 580224 656888
rect 3516 647216 3568 647222
rect 3516 647158 3568 647164
rect 67364 647216 67416 647222
rect 67364 647158 67416 647164
rect 67376 646649 67404 647158
rect 67362 646640 67418 646649
rect 67362 646575 67418 646584
rect 521028 645833 521056 656882
rect 521014 645824 521070 645833
rect 521014 645759 521070 645768
rect 3422 645144 3478 645153
rect 3422 645079 3478 645088
rect 3436 636206 3464 645079
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 520924 643136 520976 643142
rect 520924 643078 520976 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 3424 636200 3476 636206
rect 3424 636142 3476 636148
rect 67364 636200 67416 636206
rect 67364 636142 67416 636148
rect 67376 635497 67404 636142
rect 67362 635488 67418 635497
rect 67362 635423 67418 635432
rect 520936 634545 520964 643078
rect 520922 634536 520978 634545
rect 520922 634471 520978 634480
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3436 624986 3464 632023
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 520924 630692 520976 630698
rect 520924 630634 520976 630640
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 3424 624980 3476 624986
rect 3424 624922 3476 624928
rect 67364 624980 67416 624986
rect 67364 624922 67416 624928
rect 67376 624209 67404 624922
rect 67362 624200 67418 624209
rect 67362 624135 67418 624144
rect 520936 622985 520964 630634
rect 520922 622976 520978 622985
rect 520922 622911 520978 622920
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3436 614106 3464 619103
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 617030 580212 617471
rect 520280 617024 520332 617030
rect 520280 616966 520332 616972
rect 580172 617024 580224 617030
rect 580172 616966 580224 616972
rect 3424 614100 3476 614106
rect 3424 614042 3476 614048
rect 66904 614100 66956 614106
rect 66904 614042 66956 614048
rect 66916 613057 66944 614042
rect 66902 613048 66958 613057
rect 66902 612983 66958 612992
rect 520292 611697 520320 616966
rect 520278 611688 520334 611697
rect 520278 611623 520334 611632
rect 4066 606112 4122 606121
rect 4066 606047 4122 606056
rect 4080 603090 4108 606047
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 521108 603152 521160 603158
rect 521108 603094 521160 603100
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 4068 603084 4120 603090
rect 4068 603026 4120 603032
rect 66444 603084 66496 603090
rect 66444 603026 66496 603032
rect 66456 601905 66484 603026
rect 66442 601896 66498 601905
rect 66442 601831 66498 601840
rect 521120 600273 521148 603094
rect 521106 600264 521162 600273
rect 521106 600199 521162 600208
rect 3422 593056 3478 593065
rect 3422 592991 3478 593000
rect 3436 592006 3464 592991
rect 3424 592000 3476 592006
rect 3424 591942 3476 591948
rect 66996 592000 67048 592006
rect 66996 591942 67048 591948
rect 67008 590753 67036 591942
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 66994 590744 67050 590753
rect 579816 590714 579844 590951
rect 66994 590679 67050 590688
rect 521568 590708 521620 590714
rect 521568 590650 521620 590656
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 521580 588849 521608 590650
rect 521566 588840 521622 588849
rect 521566 588775 521622 588784
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 579630 3464 579935
rect 3424 579624 3476 579630
rect 67180 579624 67232 579630
rect 3424 579566 3476 579572
rect 67178 579592 67180 579601
rect 67232 579592 67234 579601
rect 67178 579527 67234 579536
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 521566 577552 521622 577561
rect 580184 577522 580212 577623
rect 521566 577487 521568 577496
rect 521620 577487 521622 577496
rect 580172 577516 580224 577522
rect 521568 577458 521620 577464
rect 580172 577458 580224 577464
rect 67362 568304 67418 568313
rect 67362 568239 67418 568248
rect 67376 567254 67404 568239
rect 4068 567248 4120 567254
rect 4068 567190 4120 567196
rect 67364 567248 67416 567254
rect 67364 567190 67416 567196
rect 4080 566953 4108 567190
rect 4066 566944 4122 566953
rect 4066 566879 4122 566888
rect 520738 566128 520794 566137
rect 520738 566063 520794 566072
rect 520752 564398 520780 566063
rect 520740 564392 520792 564398
rect 580172 564392 580224 564398
rect 520740 564334 520792 564340
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 67362 557288 67418 557297
rect 67362 557223 67418 557232
rect 67376 556238 67404 557223
rect 3424 556232 3476 556238
rect 3424 556174 3476 556180
rect 67364 556232 67416 556238
rect 67364 556174 67416 556180
rect 3436 553897 3464 556174
rect 521014 554704 521070 554713
rect 521014 554639 521070 554648
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 521028 552022 521056 554639
rect 521016 552016 521068 552022
rect 521016 551958 521068 551964
rect 579988 552016 580040 552022
rect 579988 551958 580040 551964
rect 580000 551177 580028 551958
rect 579986 551168 580042 551177
rect 579986 551103 580042 551112
rect 66626 546000 66682 546009
rect 66626 545935 66682 545944
rect 66640 545222 66668 545935
rect 2964 545216 3016 545222
rect 2964 545158 3016 545164
rect 66628 545216 66680 545222
rect 66628 545158 66680 545164
rect 2976 540841 3004 545158
rect 520922 543280 520978 543289
rect 520922 543215 520978 543224
rect 2962 540832 3018 540841
rect 2962 540767 3018 540776
rect 520936 538218 520964 543215
rect 520924 538212 520976 538218
rect 520924 538154 520976 538160
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 67362 534848 67418 534857
rect 67362 534783 67418 534792
rect 67376 534138 67404 534783
rect 3424 534132 3476 534138
rect 3424 534074 3476 534080
rect 67364 534132 67416 534138
rect 67364 534074 67416 534080
rect 3436 527921 3464 534074
rect 520922 531992 520978 532001
rect 520922 531927 520978 531936
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 520936 525774 520964 531927
rect 520924 525768 520976 525774
rect 520924 525710 520976 525716
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 66442 523696 66498 523705
rect 66442 523631 66498 523640
rect 66456 523054 66484 523631
rect 3424 523048 3476 523054
rect 3424 522990 3476 522996
rect 66444 523048 66496 523054
rect 66444 522990 66496 522996
rect 3436 514865 3464 522990
rect 520922 520568 520978 520577
rect 520922 520503 520978 520512
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 67362 512408 67418 512417
rect 67362 512343 67418 512352
rect 67376 512038 67404 512343
rect 3424 512032 3476 512038
rect 3424 511974 3476 511980
rect 67364 512032 67416 512038
rect 67364 511974 67416 511980
rect 3436 501809 3464 511974
rect 520936 511834 520964 520503
rect 520924 511828 520976 511834
rect 520924 511770 520976 511776
rect 580172 511828 580224 511834
rect 580172 511770 580224 511776
rect 580184 511329 580212 511770
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 521014 509144 521070 509153
rect 521014 509079 521070 509088
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 67454 501392 67510 501401
rect 67454 501327 67510 501336
rect 67468 501158 67496 501327
rect 3516 501152 3568 501158
rect 3516 501094 3568 501100
rect 67456 501152 67508 501158
rect 67456 501094 67508 501100
rect 3424 489932 3476 489938
rect 3424 489874 3476 489880
rect 3436 475697 3464 489874
rect 3528 488753 3556 501094
rect 521028 498166 521056 509079
rect 521016 498160 521068 498166
rect 521016 498102 521068 498108
rect 580172 498160 580224 498166
rect 580172 498102 580224 498108
rect 580184 498001 580212 498102
rect 580170 497992 580226 498001
rect 580170 497927 580226 497936
rect 520922 497856 520978 497865
rect 520922 497791 520978 497800
rect 67454 490104 67510 490113
rect 67454 490039 67510 490048
rect 67468 489938 67496 490039
rect 67456 489932 67508 489938
rect 67456 489874 67508 489880
rect 3514 488744 3570 488753
rect 3514 488679 3570 488688
rect 520936 485722 520964 497791
rect 521014 486296 521070 486305
rect 521014 486231 521070 486240
rect 520924 485716 520976 485722
rect 520924 485658 520976 485664
rect 67362 479088 67418 479097
rect 67362 479023 67418 479032
rect 67376 478922 67404 479023
rect 3516 478916 3568 478922
rect 3516 478858 3568 478864
rect 67364 478916 67416 478922
rect 67364 478858 67416 478864
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3424 466472 3476 466478
rect 3424 466414 3476 466420
rect 3436 449585 3464 466414
rect 3528 462641 3556 478858
rect 520922 475008 520978 475017
rect 520922 474943 520978 474952
rect 66994 467800 67050 467809
rect 66994 467735 67050 467744
rect 67008 466478 67036 467735
rect 66996 466472 67048 466478
rect 66996 466414 67048 466420
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 520936 458182 520964 474943
rect 521028 471986 521056 486231
rect 580172 485716 580224 485722
rect 580172 485658 580224 485664
rect 580184 484673 580212 485658
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 521016 471980 521068 471986
rect 521016 471922 521068 471928
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 521106 463584 521162 463593
rect 521106 463519 521162 463528
rect 520924 458176 520976 458182
rect 520924 458118 520976 458124
rect 67362 456648 67418 456657
rect 67362 456583 67418 456592
rect 67376 455462 67404 456583
rect 3516 455456 3568 455462
rect 3516 455398 3568 455404
rect 67364 455456 67416 455462
rect 67364 455398 67416 455404
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3424 444576 3476 444582
rect 3424 444518 3476 444524
rect 3436 423609 3464 444518
rect 3528 436665 3556 455398
rect 521014 452160 521070 452169
rect 521014 452095 521070 452104
rect 66718 445496 66774 445505
rect 66718 445431 66774 445440
rect 66732 444582 66760 445431
rect 66720 444576 66772 444582
rect 66720 444518 66772 444524
rect 520922 440872 520978 440881
rect 520922 440807 520978 440816
rect 3514 436656 3570 436665
rect 3514 436591 3570 436600
rect 67178 434344 67234 434353
rect 67178 434279 67234 434288
rect 67192 433362 67220 434279
rect 3608 433356 3660 433362
rect 3608 433298 3660 433304
rect 67180 433356 67232 433362
rect 67180 433298 67232 433304
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3424 411392 3476 411398
rect 3424 411334 3476 411340
rect 3436 384441 3464 411334
rect 3528 397497 3556 422282
rect 3620 410553 3648 433298
rect 66810 423192 66866 423201
rect 66810 423127 66866 423136
rect 66824 422346 66852 423127
rect 66812 422340 66864 422346
rect 66812 422282 66864 422288
rect 520936 419354 520964 440807
rect 521028 431866 521056 452095
rect 521120 445738 521148 463519
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 521108 445732 521160 445738
rect 521108 445674 521160 445680
rect 580172 445732 580224 445738
rect 580172 445674 580224 445680
rect 580184 444825 580212 445674
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 521016 431860 521068 431866
rect 521016 431802 521068 431808
rect 580172 431860 580224 431866
rect 580172 431802 580224 431808
rect 580184 431633 580212 431802
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 521014 429448 521070 429457
rect 521014 429383 521070 429392
rect 520924 419348 520976 419354
rect 520924 419290 520976 419296
rect 520922 418160 520978 418169
rect 520922 418095 520978 418104
rect 67270 411904 67326 411913
rect 67270 411839 67326 411848
rect 67284 411398 67312 411839
rect 67272 411392 67324 411398
rect 67272 411334 67324 411340
rect 3606 410544 3662 410553
rect 3606 410479 3662 410488
rect 67454 400888 67510 400897
rect 67454 400823 67510 400832
rect 67468 400246 67496 400823
rect 3608 400240 3660 400246
rect 3608 400182 3660 400188
rect 67456 400240 67508 400246
rect 67456 400182 67508 400188
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3516 389224 3568 389230
rect 3516 389166 3568 389172
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3424 378208 3476 378214
rect 3424 378150 3476 378156
rect 3436 345409 3464 378150
rect 3528 358465 3556 389166
rect 3620 371385 3648 400182
rect 520936 391950 520964 418095
rect 521028 405686 521056 429383
rect 580172 419348 580224 419354
rect 580172 419290 580224 419296
rect 580184 418305 580212 419290
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 521106 406736 521162 406745
rect 521106 406671 521162 406680
rect 521016 405680 521068 405686
rect 521016 405622 521068 405628
rect 521014 395312 521070 395321
rect 521014 395247 521070 395256
rect 520924 391944 520976 391950
rect 520924 391886 520976 391892
rect 67362 389600 67418 389609
rect 67362 389535 67418 389544
rect 67376 389230 67404 389535
rect 67364 389224 67416 389230
rect 67364 389166 67416 389172
rect 520922 384024 520978 384033
rect 520922 383959 520978 383968
rect 67362 378448 67418 378457
rect 67362 378383 67418 378392
rect 67376 378214 67404 378383
rect 67364 378208 67416 378214
rect 67364 378150 67416 378156
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 67362 367296 67418 367305
rect 67362 367231 67418 367240
rect 67376 367130 67404 367231
rect 3700 367124 3752 367130
rect 3700 367066 3752 367072
rect 67364 367124 67416 367130
rect 67364 367066 67416 367072
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3608 356108 3660 356114
rect 3608 356050 3660 356056
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3516 343664 3568 343670
rect 3516 343606 3568 343612
rect 3424 332648 3476 332654
rect 3424 332590 3476 332596
rect 3436 293185 3464 332590
rect 3528 306241 3556 343606
rect 3620 319297 3648 356050
rect 3712 332353 3740 367066
rect 67362 356144 67418 356153
rect 67362 356079 67364 356088
rect 67416 356079 67418 356088
rect 67364 356050 67416 356056
rect 520936 353258 520964 383959
rect 521028 365702 521056 395247
rect 521120 379506 521148 406671
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 391944 580224 391950
rect 580172 391886 580224 391892
rect 580184 391785 580212 391886
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 521108 379500 521160 379506
rect 521108 379442 521160 379448
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 521198 372464 521254 372473
rect 521198 372399 521254 372408
rect 521016 365696 521068 365702
rect 521016 365638 521068 365644
rect 521106 361176 521162 361185
rect 521106 361111 521162 361120
rect 520924 353252 520976 353258
rect 520924 353194 520976 353200
rect 521014 349888 521070 349897
rect 521014 349823 521070 349832
rect 67362 344992 67418 345001
rect 67362 344927 67418 344936
rect 67376 343670 67404 344927
rect 67364 343664 67416 343670
rect 67364 343606 67416 343612
rect 520922 338328 520978 338337
rect 520922 338263 520978 338272
rect 67178 333840 67234 333849
rect 67178 333775 67234 333784
rect 67192 332654 67220 333775
rect 67180 332648 67232 332654
rect 67180 332590 67232 332596
rect 3698 332344 3754 332353
rect 3698 332279 3754 332288
rect 67362 322688 67418 322697
rect 67362 322623 67418 322632
rect 67376 321638 67404 322623
rect 3700 321632 3752 321638
rect 3700 321574 3752 321580
rect 67364 321632 67416 321638
rect 67364 321574 67416 321580
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3608 310548 3660 310554
rect 3608 310490 3660 310496
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 299532 3568 299538
rect 3516 299474 3568 299480
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3424 288448 3476 288454
rect 3424 288390 3476 288396
rect 3436 241097 3464 288390
rect 3528 254153 3556 299474
rect 3620 267209 3648 310490
rect 3712 280129 3740 321574
rect 66718 311400 66774 311409
rect 66718 311335 66774 311344
rect 66732 310554 66760 311335
rect 66720 310548 66772 310554
rect 66720 310490 66772 310496
rect 67362 300248 67418 300257
rect 67362 300183 67418 300192
rect 67376 299538 67404 300183
rect 67364 299532 67416 299538
rect 67364 299474 67416 299480
rect 520936 299470 520964 338263
rect 521028 313274 521056 349823
rect 521120 325650 521148 361111
rect 521212 339386 521240 372399
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 521200 339380 521252 339386
rect 521200 339322 521252 339328
rect 580172 339380 580224 339386
rect 580172 339322 580224 339328
rect 580184 338609 580212 339322
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 521198 327040 521254 327049
rect 521198 326975 521254 326984
rect 521108 325644 521160 325650
rect 521108 325586 521160 325592
rect 521106 315616 521162 315625
rect 521106 315551 521162 315560
rect 521016 313268 521068 313274
rect 521016 313210 521068 313216
rect 521014 304192 521070 304201
rect 521014 304127 521070 304136
rect 520924 299464 520976 299470
rect 520924 299406 520976 299412
rect 520922 292904 520978 292913
rect 520922 292839 520978 292848
rect 66442 289096 66498 289105
rect 66442 289031 66498 289040
rect 66456 288454 66484 289031
rect 66444 288448 66496 288454
rect 66444 288390 66496 288396
rect 3698 280120 3754 280129
rect 3698 280055 3754 280064
rect 67362 277944 67418 277953
rect 67362 277879 67418 277888
rect 67376 277574 67404 277879
rect 3792 277568 3844 277574
rect 3792 277510 3844 277516
rect 67364 277568 67416 277574
rect 67364 277510 67416 277516
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3700 266416 3752 266422
rect 3700 266358 3752 266364
rect 3608 255332 3660 255338
rect 3608 255274 3660 255280
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 244384 3568 244390
rect 3516 244326 3568 244332
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3424 233300 3476 233306
rect 3424 233242 3476 233248
rect 3436 175953 3464 233242
rect 3528 188873 3556 244326
rect 3620 201929 3648 255274
rect 3712 214985 3740 266358
rect 3804 228041 3832 277510
rect 67362 266792 67418 266801
rect 67362 266727 67418 266736
rect 67376 266422 67404 266727
rect 67364 266416 67416 266422
rect 67364 266358 67416 266364
rect 67362 255640 67418 255649
rect 67362 255575 67418 255584
rect 67376 255338 67404 255575
rect 67364 255332 67416 255338
rect 67364 255274 67416 255280
rect 520936 245614 520964 292839
rect 521028 259418 521056 304127
rect 521120 273222 521148 315551
rect 521212 285530 521240 326975
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 521200 285524 521252 285530
rect 521200 285466 521252 285472
rect 580172 285524 580224 285530
rect 580172 285466 580224 285472
rect 580184 285433 580212 285466
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 521290 281480 521346 281489
rect 521290 281415 521346 281424
rect 521108 273216 521160 273222
rect 521108 273158 521160 273164
rect 521198 270056 521254 270065
rect 521198 269991 521254 270000
rect 521016 259412 521068 259418
rect 521016 259354 521068 259360
rect 521106 258768 521162 258777
rect 521106 258703 521162 258712
rect 521014 247344 521070 247353
rect 521014 247279 521070 247288
rect 520924 245608 520976 245614
rect 520924 245550 520976 245556
rect 67362 244488 67418 244497
rect 67362 244423 67418 244432
rect 67376 244390 67404 244423
rect 67364 244384 67416 244390
rect 67364 244326 67416 244332
rect 520922 235920 520978 235929
rect 520922 235855 520978 235864
rect 67178 233336 67234 233345
rect 67178 233271 67180 233280
rect 67232 233271 67234 233280
rect 67180 233242 67232 233248
rect 3790 228032 3846 228041
rect 3790 227967 3846 227976
rect 67362 222048 67418 222057
rect 67362 221983 67418 221992
rect 67376 220998 67404 221983
rect 3884 220992 3936 220998
rect 3884 220934 3936 220940
rect 67364 220992 67416 220998
rect 67364 220934 67416 220940
rect 3698 214976 3754 214985
rect 3698 214911 3754 214920
rect 3792 209840 3844 209846
rect 3792 209782 3844 209788
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3700 198756 3752 198762
rect 3700 198698 3752 198704
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3608 187808 3660 187814
rect 3608 187750 3660 187756
rect 3516 176724 3568 176730
rect 3516 176666 3568 176672
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 3424 165640 3476 165646
rect 3424 165582 3476 165588
rect 3436 97617 3464 165582
rect 3528 110673 3556 176666
rect 3620 123729 3648 187750
rect 3712 136785 3740 198698
rect 3804 149841 3832 209782
rect 3896 162897 3924 220934
rect 67362 210896 67418 210905
rect 67362 210831 67418 210840
rect 67376 209846 67404 210831
rect 67364 209840 67416 209846
rect 67364 209782 67416 209788
rect 67362 199744 67418 199753
rect 67362 199679 67418 199688
rect 67376 198762 67404 199679
rect 67364 198756 67416 198762
rect 67364 198698 67416 198704
rect 67454 188592 67510 188601
rect 67454 188527 67510 188536
rect 67468 187814 67496 188527
rect 67456 187808 67508 187814
rect 67456 187750 67508 187756
rect 520936 179382 520964 235855
rect 521028 193050 521056 247279
rect 521120 206990 521148 258703
rect 521212 219434 521240 269991
rect 521304 233238 521332 281415
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 521292 233232 521344 233238
rect 521292 233174 521344 233180
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 521382 224496 521438 224505
rect 521382 224431 521438 224440
rect 521200 219428 521252 219434
rect 521200 219370 521252 219376
rect 521290 213208 521346 213217
rect 521290 213143 521346 213152
rect 521108 206984 521160 206990
rect 521108 206926 521160 206932
rect 521198 201784 521254 201793
rect 521198 201719 521254 201728
rect 521016 193044 521068 193050
rect 521016 192986 521068 192992
rect 521106 190360 521162 190369
rect 521106 190295 521162 190304
rect 520924 179376 520976 179382
rect 520924 179318 520976 179324
rect 521014 179072 521070 179081
rect 521014 179007 521070 179016
rect 67362 177440 67418 177449
rect 67362 177375 67418 177384
rect 67376 176730 67404 177375
rect 67364 176724 67416 176730
rect 67364 176666 67416 176672
rect 520922 167648 520978 167657
rect 520922 167583 520978 167592
rect 67362 166288 67418 166297
rect 67362 166223 67418 166232
rect 67376 165646 67404 166223
rect 67364 165640 67416 165646
rect 67364 165582 67416 165588
rect 3882 162888 3938 162897
rect 3882 162823 3938 162832
rect 67270 155136 67326 155145
rect 67270 155071 67326 155080
rect 67284 154630 67312 155071
rect 3976 154624 4028 154630
rect 3976 154566 4028 154572
rect 67272 154624 67324 154630
rect 67272 154566 67324 154572
rect 3790 149832 3846 149841
rect 3790 149767 3846 149776
rect 3884 143744 3936 143750
rect 3884 143686 3936 143692
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 3792 132524 3844 132530
rect 3792 132466 3844 132472
rect 3606 123720 3662 123729
rect 3606 123655 3662 123664
rect 3700 121508 3752 121514
rect 3700 121450 3752 121456
rect 3514 110664 3570 110673
rect 3514 110599 3570 110608
rect 3608 109064 3660 109070
rect 3608 109006 3660 109012
rect 3516 98048 3568 98054
rect 3516 97990 3568 97996
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3424 88392 3476 88398
rect 3424 88334 3476 88340
rect 3436 6497 3464 88334
rect 3528 19417 3556 97990
rect 3620 32473 3648 109006
rect 3712 45529 3740 121450
rect 3804 58585 3832 132466
rect 3896 71641 3924 143686
rect 3988 84697 4016 154566
rect 67362 143848 67418 143857
rect 67362 143783 67418 143792
rect 67376 143750 67404 143783
rect 67364 143744 67416 143750
rect 67364 143686 67416 143692
rect 67178 132832 67234 132841
rect 67178 132767 67234 132776
rect 67192 132530 67220 132767
rect 67180 132524 67232 132530
rect 67180 132466 67232 132472
rect 67362 121544 67418 121553
rect 67362 121479 67364 121488
rect 67416 121479 67418 121488
rect 67364 121450 67416 121456
rect 67362 110392 67418 110401
rect 67362 110327 67418 110336
rect 67376 109070 67404 110327
rect 67364 109064 67416 109070
rect 67364 109006 67416 109012
rect 520936 100570 520964 167583
rect 521028 113082 521056 179007
rect 521120 126954 521148 190295
rect 521212 139398 521240 201719
rect 521304 153202 521332 213143
rect 521396 166938 521424 224431
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193044 580224 193050
rect 580172 192986 580224 192992
rect 580184 192545 580212 192986
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 521384 166932 521436 166938
rect 521384 166874 521436 166880
rect 580172 166932 580224 166938
rect 580172 166874 580224 166880
rect 580184 165889 580212 166874
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 521474 156224 521530 156233
rect 521474 156159 521530 156168
rect 521292 153196 521344 153202
rect 521292 153138 521344 153144
rect 521382 144800 521438 144809
rect 521382 144735 521438 144744
rect 521200 139392 521252 139398
rect 521200 139334 521252 139340
rect 521290 133512 521346 133521
rect 521290 133447 521346 133456
rect 521108 126948 521160 126954
rect 521108 126890 521160 126896
rect 521198 122088 521254 122097
rect 521198 122023 521254 122032
rect 521016 113076 521068 113082
rect 521016 113018 521068 113024
rect 521106 110664 521162 110673
rect 521106 110599 521162 110608
rect 520924 100564 520976 100570
rect 520924 100506 520976 100512
rect 521014 99376 521070 99385
rect 521014 99311 521070 99320
rect 67178 99240 67234 99249
rect 67178 99175 67234 99184
rect 67192 98054 67220 99175
rect 67180 98048 67232 98054
rect 67180 97990 67232 97996
rect 67454 89176 67510 89185
rect 67454 89111 67510 89120
rect 67468 88398 67496 89111
rect 520922 88904 520978 88913
rect 520922 88839 520978 88848
rect 67456 88392 67508 88398
rect 67456 88334 67508 88340
rect 70860 87938 70888 88049
rect 70780 87910 70888 87938
rect 70780 87802 70808 87910
rect 70952 87802 70980 88049
rect 70412 87774 70808 87802
rect 70872 87774 70980 87802
rect 71780 87802 71808 88049
rect 72700 87802 72728 88049
rect 71780 87774 71820 87802
rect 18604 85128 18656 85134
rect 18604 85070 18656 85076
rect 7564 84992 7616 84998
rect 7564 84934 7616 84940
rect 3974 84688 4030 84697
rect 3974 84623 4030 84632
rect 3882 71632 3938 71641
rect 3882 71567 3938 71576
rect 3790 58576 3846 58585
rect 3790 58511 3846 58520
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 572 5024 624 5030
rect 572 4966 624 4972
rect 584 480 612 4966
rect 1688 480 1716 5102
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2884 480 2912 5034
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 480 4108 4762
rect 7576 4146 7604 84934
rect 10324 83496 10376 83502
rect 10324 83438 10376 83444
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 4082
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 480 7696 3402
rect 8772 480 8800 3538
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9968 480 9996 3470
rect 10336 3466 10364 83438
rect 14464 80708 14516 80714
rect 14464 80650 14516 80656
rect 12348 77988 12400 77994
rect 12348 77930 12400 77936
rect 10968 57248 11020 57254
rect 10968 57190 11020 57196
rect 10980 3534 11008 57190
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11150 3496 11206 3505
rect 10324 3460 10376 3466
rect 11150 3431 11206 3440
rect 10324 3402 10376 3408
rect 11164 480 11192 3431
rect 12360 480 12388 77930
rect 14476 3602 14504 80650
rect 15844 68332 15896 68338
rect 15844 68274 15896 68280
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13556 480 13584 2994
rect 14752 480 14780 4014
rect 15856 3058 15884 68274
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 480 15976 3538
rect 17880 3126 17908 17206
rect 18616 4078 18644 85070
rect 19984 85060 20036 85066
rect 19984 85002 20036 85008
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 19260 3534 19288 29582
rect 19996 3602 20024 85002
rect 62028 83564 62080 83570
rect 62028 83506 62080 83512
rect 59268 80776 59320 80782
rect 59268 80718 59320 80724
rect 30288 75268 30340 75274
rect 30288 75210 30340 75216
rect 28908 65544 28960 65550
rect 28908 65486 28960 65492
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 20626 3632 20682 3641
rect 19984 3596 20036 3602
rect 20626 3567 20682 3576
rect 19984 3538 20036 3544
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17052 480 17080 3062
rect 18248 480 18276 3470
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 480 19472 3402
rect 20640 480 20668 3567
rect 21836 480 21864 8910
rect 23400 6914 23428 32370
rect 23032 6886 23428 6914
rect 23032 480 23060 6886
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 25318 3768 25374 3777
rect 25318 3703 25374 3712
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3703
rect 26528 480 26556 6122
rect 28920 3602 28948 65486
rect 30300 6914 30328 75210
rect 34428 73840 34480 73846
rect 34428 73782 34480 73788
rect 32404 62824 32456 62830
rect 32404 62766 32456 62772
rect 30116 6886 30328 6914
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27724 480 27752 3538
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30116 480 30144 6886
rect 32416 3602 32444 62766
rect 32496 3664 32548 3670
rect 32496 3606 32548 3612
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 31312 480 31340 3538
rect 32508 1850 32536 3606
rect 34440 3602 34468 73782
rect 37188 71052 37240 71058
rect 37188 70994 37240 71000
rect 35808 37936 35860 37942
rect 35808 37878 35860 37884
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 32416 1822 32536 1850
rect 32416 480 32444 1822
rect 33612 480 33640 3538
rect 35820 3398 35848 37878
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3674
rect 37200 480 37228 70994
rect 38568 60036 38620 60042
rect 38568 59978 38620 59984
rect 38580 6914 38608 59978
rect 50988 55888 51040 55894
rect 50988 55830 51040 55836
rect 45468 35216 45520 35222
rect 45468 35158 45520 35164
rect 42708 26920 42760 26926
rect 42708 26862 42760 26868
rect 41328 14476 41380 14482
rect 41328 14418 41380 14424
rect 38396 6886 38608 6914
rect 38396 480 38424 6886
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39592 480 39620 3878
rect 41340 3398 41368 14418
rect 42720 3398 42748 26862
rect 45376 18624 45428 18630
rect 45376 18566 45428 18572
rect 43076 4004 43128 4010
rect 43076 3946 43128 3952
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3334
rect 43088 480 43116 3946
rect 45388 3398 45416 18566
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 44284 480 44312 3334
rect 45480 480 45508 35158
rect 48964 5228 49016 5234
rect 48964 5170 49016 5176
rect 47860 4752 47912 4758
rect 47860 4694 47912 4700
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 46676 480 46704 4014
rect 47872 480 47900 4694
rect 48976 480 49004 5170
rect 51000 3398 51028 55830
rect 57888 53100 57940 53106
rect 57888 53042 57940 53048
rect 53748 42084 53800 42090
rect 53748 42026 53800 42032
rect 53656 21412 53708 21418
rect 53656 21354 53708 21360
rect 51356 4684 51408 4690
rect 51356 4626 51408 4632
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50172 480 50200 3334
rect 51368 480 51396 4626
rect 53668 3398 53696 21354
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 53656 3392 53708 3398
rect 53656 3334 53708 3340
rect 52564 480 52592 3334
rect 53760 480 53788 42026
rect 56048 5296 56100 5302
rect 56048 5238 56100 5244
rect 54944 4616 54996 4622
rect 54944 4558 54996 4564
rect 54956 480 54984 4558
rect 56060 480 56088 5238
rect 57900 3398 57928 53042
rect 59280 3398 59308 80718
rect 61936 47592 61988 47598
rect 61936 47534 61988 47540
rect 60648 11756 60700 11762
rect 60648 11698 60700 11704
rect 60660 3398 60688 11698
rect 61948 3398 61976 47534
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 61936 3392 61988 3398
rect 61936 3334 61988 3340
rect 57256 480 57284 3334
rect 58452 480 58480 3334
rect 59648 480 59676 3334
rect 60844 480 60872 3334
rect 62040 480 62068 83506
rect 70216 78056 70268 78062
rect 70216 77998 70268 78004
rect 64788 50380 64840 50386
rect 64788 50322 64840 50328
rect 63224 5364 63276 5370
rect 63224 5306 63276 5312
rect 63236 480 63264 5306
rect 64800 3398 64828 50322
rect 68928 44872 68980 44878
rect 68928 44814 68980 44820
rect 66720 9036 66772 9042
rect 66720 8978 66772 8984
rect 65524 4548 65576 4554
rect 65524 4490 65576 4496
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64340 480 64368 3334
rect 65536 480 65564 4490
rect 66732 480 66760 8978
rect 68940 3398 68968 44814
rect 70228 16574 70256 77998
rect 70228 16546 70348 16574
rect 69112 4480 69164 4486
rect 69112 4422 69164 4428
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 67928 480 67956 3334
rect 69124 480 69152 4422
rect 70320 480 70348 16546
rect 70412 5166 70440 87774
rect 70872 84194 70900 87774
rect 70504 84166 70900 84194
rect 70400 5160 70452 5166
rect 70400 5102 70452 5108
rect 70504 5030 70532 84166
rect 71688 39364 71740 39370
rect 71688 39306 71740 39312
rect 71700 6914 71728 39306
rect 71516 6886 71728 6914
rect 70492 5024 70544 5030
rect 70492 4966 70544 4972
rect 71516 480 71544 6886
rect 71792 5098 71820 87774
rect 72620 87774 72728 87802
rect 73160 87848 73212 87854
rect 73620 87802 73648 88049
rect 74448 87854 74476 88049
rect 73160 87790 73212 87796
rect 72620 84194 72648 87774
rect 71884 84166 72648 84194
rect 71884 83502 71912 84166
rect 71872 83496 71924 83502
rect 71872 83438 71924 83444
rect 73172 17270 73200 87790
rect 73540 87774 73648 87802
rect 74436 87848 74488 87854
rect 75368 87802 75396 88049
rect 76288 87802 76316 88049
rect 74436 87790 74488 87796
rect 75288 87774 75396 87802
rect 76208 87774 76316 87802
rect 77208 87802 77236 88049
rect 78128 87802 78156 88049
rect 78680 87848 78732 87854
rect 77208 87774 77248 87802
rect 78128 87774 78168 87802
rect 79048 87802 79076 88049
rect 79968 87854 79996 88049
rect 78680 87790 78732 87796
rect 73540 84194 73568 87774
rect 75288 84194 75316 87774
rect 76208 86954 76236 87774
rect 73264 84166 73568 84194
rect 74552 84166 75316 84194
rect 75932 86926 76236 86954
rect 73264 77994 73292 84166
rect 73252 77988 73304 77994
rect 73252 77930 73304 77936
rect 74448 17332 74500 17338
rect 74448 17274 74500 17280
rect 73160 17264 73212 17270
rect 73160 17206 73212 17212
rect 73068 11824 73120 11830
rect 73068 11766 73120 11772
rect 71780 5092 71832 5098
rect 71780 5034 71832 5040
rect 73080 3398 73108 11766
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 72620 480 72648 3334
rect 74460 2922 74488 17274
rect 74552 8974 74580 84166
rect 75828 75200 75880 75206
rect 75828 75142 75880 75148
rect 74540 8968 74592 8974
rect 74540 8910 74592 8916
rect 75840 3398 75868 75142
rect 75932 6186 75960 86926
rect 77220 86154 77248 87774
rect 76012 86148 76064 86154
rect 76012 86090 76064 86096
rect 77208 86148 77260 86154
rect 77208 86090 77260 86096
rect 76024 75274 76052 86090
rect 78140 85542 78168 87774
rect 76564 85536 76616 85542
rect 76564 85478 76616 85484
rect 78128 85536 78180 85542
rect 78128 85478 78180 85484
rect 76012 75268 76064 75274
rect 76012 75210 76064 75216
rect 76576 73846 76604 85478
rect 76564 73840 76616 73846
rect 76564 73782 76616 73788
rect 78588 17264 78640 17270
rect 78588 17206 78640 17212
rect 76196 6248 76248 6254
rect 76196 6190 76248 6196
rect 75920 6180 75972 6186
rect 75920 6122 75972 6128
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75828 3392 75880 3398
rect 75828 3334 75880 3340
rect 73804 2916 73856 2922
rect 73804 2858 73856 2864
rect 74448 2916 74500 2922
rect 74448 2858 74500 2864
rect 73816 480 73844 2858
rect 75012 480 75040 3334
rect 76208 480 76236 6190
rect 77392 6180 77444 6186
rect 77392 6122 77444 6128
rect 77404 480 77432 6122
rect 78600 480 78628 17206
rect 78692 14482 78720 87790
rect 78968 87774 79076 87802
rect 79956 87848 80008 87854
rect 79956 87790 80008 87796
rect 80888 87802 80916 88049
rect 81716 87802 81744 88049
rect 82636 87802 82664 88049
rect 83556 87802 83584 88049
rect 84476 87802 84504 88049
rect 85396 87802 85424 88049
rect 86316 87802 86344 88049
rect 87236 87802 87264 88049
rect 88156 87802 88184 88049
rect 88984 87802 89012 88049
rect 89904 87802 89932 88049
rect 90824 87802 90852 88049
rect 91744 87802 91772 88049
rect 92664 87802 92692 88049
rect 80888 87774 80928 87802
rect 78968 84194 78996 87774
rect 80900 85542 80928 87774
rect 81636 87774 81744 87802
rect 82556 87774 82664 87802
rect 83476 87774 83584 87802
rect 84396 87774 84504 87802
rect 85316 87774 85424 87802
rect 86236 87774 86344 87802
rect 86972 87774 87264 87802
rect 88076 87774 88184 87802
rect 88904 87774 89012 87802
rect 89732 87774 89932 87802
rect 90744 87774 90852 87802
rect 91664 87774 91772 87802
rect 92584 87774 92692 87802
rect 93584 87802 93612 88049
rect 94504 87802 94532 88049
rect 95424 87802 95452 88049
rect 96252 87802 96280 88049
rect 97172 87802 97200 88049
rect 98092 87802 98120 88049
rect 99012 87802 99040 88049
rect 99932 87802 99960 88049
rect 100852 87802 100880 88049
rect 101772 87802 101800 88049
rect 102692 87802 102720 88049
rect 93584 87774 93624 87802
rect 94504 87774 94544 87802
rect 95424 87774 95464 87802
rect 96252 87774 96292 87802
rect 97172 87774 97212 87802
rect 98092 87774 98132 87802
rect 99012 87774 99052 87802
rect 99932 87774 99972 87802
rect 100852 87774 100892 87802
rect 81636 86954 81664 87774
rect 81452 86926 81664 86954
rect 79324 85536 79376 85542
rect 79324 85478 79376 85484
rect 80888 85536 80940 85542
rect 80888 85478 80940 85484
rect 78784 84166 78996 84194
rect 78784 71058 78812 84166
rect 78772 71052 78824 71058
rect 78772 70994 78824 71000
rect 79336 18630 79364 85478
rect 81348 18692 81400 18698
rect 81348 18634 81400 18640
rect 79324 18624 79376 18630
rect 79324 18566 79376 18572
rect 78680 14476 78732 14482
rect 78680 14418 78732 14424
rect 79692 8968 79744 8974
rect 79692 8910 79744 8916
rect 79704 480 79732 8910
rect 81360 3398 81388 18634
rect 81452 4758 81480 86926
rect 82556 84194 82584 87774
rect 83476 84194 83504 87774
rect 84396 84266 84424 87774
rect 81544 84166 82584 84194
rect 82832 84166 83504 84194
rect 84120 84238 84424 84266
rect 81440 4752 81492 4758
rect 81440 4694 81492 4700
rect 81544 4690 81572 84166
rect 82728 18624 82780 18630
rect 82728 18566 82780 18572
rect 81532 4684 81584 4690
rect 81532 4626 81584 4632
rect 82740 3398 82768 18566
rect 82832 4622 82860 84166
rect 84120 80782 84148 84238
rect 85316 84194 85344 87774
rect 86236 84194 86264 87774
rect 84304 84166 85344 84194
rect 85592 84166 86264 84194
rect 84304 83570 84332 84166
rect 84292 83564 84344 83570
rect 84292 83506 84344 83512
rect 84108 80776 84160 80782
rect 84108 80718 84160 80724
rect 84108 14544 84160 14550
rect 84108 14486 84160 14492
rect 82820 4616 82872 4622
rect 82820 4558 82872 4564
rect 84120 3398 84148 14486
rect 85488 14476 85540 14482
rect 85488 14418 85540 14424
rect 85500 3398 85528 14418
rect 85592 4554 85620 84166
rect 86868 5568 86920 5574
rect 86868 5510 86920 5516
rect 85580 4548 85632 4554
rect 85580 4490 85632 4496
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 82084 3392 82136 3398
rect 82084 3334 82136 3340
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3334
rect 83292 480 83320 3334
rect 84488 480 84516 3334
rect 85684 480 85712 4082
rect 86880 480 86908 5510
rect 86972 4486 87000 87774
rect 88076 84194 88104 87774
rect 88904 84194 88932 87774
rect 87064 84166 88104 84194
rect 88352 84166 88932 84194
rect 87064 11830 87092 84166
rect 88248 24132 88300 24138
rect 88248 24074 88300 24080
rect 87052 11824 87104 11830
rect 87052 11766 87104 11772
rect 88260 6914 88288 24074
rect 87984 6886 88288 6914
rect 86960 4480 87012 4486
rect 86960 4422 87012 4428
rect 87984 480 88012 6886
rect 88352 6254 88380 84166
rect 89732 8974 89760 87774
rect 90744 84194 90772 87774
rect 91664 84194 91692 87774
rect 92584 84194 92612 87774
rect 89824 84166 90772 84194
rect 91112 84166 91692 84194
rect 92492 84166 92612 84194
rect 93596 84194 93624 87774
rect 94516 85542 94544 87774
rect 95436 85542 95464 87774
rect 94504 85536 94556 85542
rect 94504 85478 94556 85484
rect 95148 85536 95200 85542
rect 95148 85478 95200 85484
rect 95424 85536 95476 85542
rect 95424 85478 95476 85484
rect 93596 84166 93808 84194
rect 89824 14550 89852 84166
rect 89812 14544 89864 14550
rect 89812 14486 89864 14492
rect 91008 11688 91060 11694
rect 91008 11630 91060 11636
rect 89720 8968 89772 8974
rect 89720 8910 89772 8916
rect 88340 6248 88392 6254
rect 88340 6190 88392 6196
rect 91020 3398 91048 11630
rect 91112 5574 91140 84166
rect 92388 73840 92440 73846
rect 92388 73782 92440 73788
rect 91100 5568 91152 5574
rect 91100 5510 91152 5516
rect 92400 3398 92428 73782
rect 92492 11694 92520 84166
rect 92480 11688 92532 11694
rect 92480 11630 92532 11636
rect 93780 5658 93808 84166
rect 95056 26988 95108 26994
rect 95056 26930 95108 26936
rect 93780 5630 93992 5658
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 92388 3392 92440 3398
rect 92388 3334 92440 3340
rect 89168 3188 89220 3194
rect 89168 3130 89220 3136
rect 89180 480 89208 3130
rect 90376 480 90404 3334
rect 91572 480 91600 3334
rect 92756 3188 92808 3194
rect 92756 3130 92808 3136
rect 92768 480 92796 3130
rect 93964 480 93992 5630
rect 95068 3482 95096 26930
rect 95160 4214 95188 85478
rect 96264 84194 96292 87774
rect 97184 85542 97212 87774
rect 98104 85542 98132 87774
rect 96436 85536 96488 85542
rect 96436 85478 96488 85484
rect 97172 85536 97224 85542
rect 97172 85478 97224 85484
rect 97908 85536 97960 85542
rect 97908 85478 97960 85484
rect 98092 85536 98144 85542
rect 98092 85478 98144 85484
rect 96264 84166 96384 84194
rect 96356 6914 96384 84166
rect 96172 6886 96384 6914
rect 96172 4690 96200 6886
rect 96160 4684 96212 4690
rect 96160 4626 96212 4632
rect 96448 4282 96476 85478
rect 96528 85196 96580 85202
rect 96528 85138 96580 85144
rect 96436 4276 96488 4282
rect 96436 4218 96488 4224
rect 95148 4208 95200 4214
rect 95148 4150 95200 4156
rect 96540 3482 96568 85138
rect 97920 5166 97948 85478
rect 99024 84194 99052 87774
rect 99944 85542 99972 87774
rect 100864 85542 100892 87774
rect 101692 87774 101800 87802
rect 102612 87774 102720 87802
rect 103520 87802 103548 88049
rect 104440 87802 104468 88049
rect 105360 87802 105388 88049
rect 103520 87774 103652 87802
rect 104440 87774 104480 87802
rect 99288 85536 99340 85542
rect 99288 85478 99340 85484
rect 99932 85536 99984 85542
rect 99932 85478 99984 85484
rect 100668 85536 100720 85542
rect 100668 85478 100720 85484
rect 100852 85536 100904 85542
rect 100852 85478 100904 85484
rect 99024 84166 99236 84194
rect 98644 6248 98696 6254
rect 98644 6190 98696 6196
rect 97908 5160 97960 5166
rect 97908 5102 97960 5108
rect 97448 4208 97500 4214
rect 97448 4150 97500 4156
rect 95068 3454 95188 3482
rect 95160 480 95188 3454
rect 96264 3454 96568 3482
rect 96264 480 96292 3454
rect 97460 480 97488 4150
rect 98656 480 98684 6190
rect 99208 5098 99236 84166
rect 99196 5092 99248 5098
rect 99196 5034 99248 5040
rect 99300 4758 99328 85478
rect 100680 5030 100708 85478
rect 101692 84194 101720 87774
rect 102048 85536 102100 85542
rect 102048 85478 102100 85484
rect 100772 84166 101720 84194
rect 100668 5024 100720 5030
rect 100668 4966 100720 4972
rect 100772 4826 100800 84166
rect 102060 4826 102088 85478
rect 102612 84194 102640 87774
rect 103520 86148 103572 86154
rect 103520 86090 103572 86096
rect 102152 84166 102640 84194
rect 102152 80714 102180 84166
rect 102140 80708 102192 80714
rect 102140 80650 102192 80656
rect 103532 29646 103560 86090
rect 103624 68338 103652 87774
rect 104452 86154 104480 87774
rect 105280 87774 105388 87802
rect 106280 87802 106308 88049
rect 107200 87802 107228 88049
rect 108120 87802 108148 88049
rect 106280 87774 106412 87802
rect 107200 87774 107240 87802
rect 104440 86148 104492 86154
rect 104440 86090 104492 86096
rect 105280 84194 105308 87774
rect 106280 86148 106332 86154
rect 106280 86090 106332 86096
rect 104912 84166 105308 84194
rect 103612 68332 103664 68338
rect 103612 68274 103664 68280
rect 104912 32434 104940 84166
rect 106292 62830 106320 86090
rect 106384 65550 106412 87774
rect 107212 86154 107240 87774
rect 108040 87774 108148 87802
rect 109040 87802 109068 88049
rect 109960 87802 109988 88049
rect 110420 87848 110472 87854
rect 109040 87774 109172 87802
rect 109960 87774 110000 87802
rect 110788 87802 110816 88049
rect 111708 87854 111736 88049
rect 112628 87938 112656 88049
rect 112364 87910 112656 87938
rect 110420 87790 110472 87796
rect 107200 86148 107252 86154
rect 107200 86090 107252 86096
rect 107568 85264 107620 85270
rect 107568 85206 107620 85212
rect 106372 65544 106424 65550
rect 106372 65486 106424 65492
rect 106280 62824 106332 62830
rect 106280 62766 106332 62772
rect 104900 32428 104952 32434
rect 104900 32370 104952 32376
rect 103520 29640 103572 29646
rect 103520 29582 103572 29588
rect 106188 11824 106240 11830
rect 106188 11766 106240 11772
rect 102232 8968 102284 8974
rect 102232 8910 102284 8916
rect 100760 4820 100812 4826
rect 100760 4762 100812 4768
rect 102048 4820 102100 4826
rect 102048 4762 102100 4768
rect 99288 4752 99340 4758
rect 99288 4694 99340 4700
rect 101036 4276 101088 4282
rect 101036 4218 101088 4224
rect 99840 3120 99892 3126
rect 99840 3062 99892 3068
rect 99852 480 99880 3062
rect 101048 480 101076 4218
rect 102244 480 102272 8910
rect 104532 4684 104584 4690
rect 104532 4626 104584 4632
rect 103336 3052 103388 3058
rect 103336 2994 103388 3000
rect 103348 480 103376 2994
rect 104544 480 104572 4626
rect 106200 2990 106228 11766
rect 107580 2990 107608 85206
rect 108040 84194 108068 87774
rect 109040 86148 109092 86154
rect 109040 86090 109092 86096
rect 107672 84166 108068 84194
rect 107672 37942 107700 84166
rect 107660 37936 107712 37942
rect 107660 37878 107712 37884
rect 109052 26926 109080 86090
rect 109144 60042 109172 87774
rect 109972 86154 110000 87774
rect 109960 86148 110012 86154
rect 109960 86090 110012 86096
rect 109132 60036 109184 60042
rect 109132 59978 109184 59984
rect 109040 26920 109092 26926
rect 109040 26862 109092 26868
rect 110328 21480 110380 21486
rect 110328 21422 110380 21428
rect 108120 5160 108172 5166
rect 108120 5102 108172 5108
rect 105728 2984 105780 2990
rect 105728 2926 105780 2932
rect 106188 2984 106240 2990
rect 106188 2926 106240 2932
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 107568 2984 107620 2990
rect 107568 2926 107620 2932
rect 105740 480 105768 2926
rect 106936 480 106964 2926
rect 108132 480 108160 5102
rect 110340 2990 110368 21422
rect 110432 5234 110460 87790
rect 110708 87774 110816 87802
rect 111696 87848 111748 87854
rect 111696 87790 111748 87796
rect 110708 84194 110736 87774
rect 112364 84194 112392 87910
rect 113548 87802 113576 88049
rect 113468 87774 113576 87802
rect 114468 87802 114496 88049
rect 115388 87938 115416 88049
rect 115124 87910 115416 87938
rect 114468 87774 114508 87802
rect 110524 84166 110736 84194
rect 111812 84166 112392 84194
rect 112444 84244 112496 84250
rect 113468 84194 113496 87774
rect 114480 84250 114508 87774
rect 112444 84186 112496 84192
rect 110524 35222 110552 84166
rect 110512 35216 110564 35222
rect 110512 35158 110564 35164
rect 111812 21418 111840 84166
rect 111800 21412 111852 21418
rect 111800 21354 111852 21360
rect 112456 11762 112484 84186
rect 113284 84166 113496 84194
rect 114468 84244 114520 84250
rect 115124 84194 115152 87910
rect 116032 87848 116084 87854
rect 116032 87790 116084 87796
rect 116308 87802 116336 88049
rect 117228 87854 117256 88049
rect 117216 87848 117268 87854
rect 115204 85536 115256 85542
rect 115204 85478 115256 85484
rect 114468 84186 114520 84192
rect 114572 84166 115152 84194
rect 113088 29640 113140 29646
rect 113088 29582 113140 29588
rect 112444 11756 112496 11762
rect 112444 11698 112496 11704
rect 113100 6914 113128 29582
rect 112824 6886 113128 6914
rect 110420 5228 110472 5234
rect 110420 5170 110472 5176
rect 111616 4752 111668 4758
rect 111616 4694 111668 4700
rect 109316 2984 109368 2990
rect 109316 2926 109368 2932
rect 110328 2984 110380 2990
rect 110328 2926 110380 2932
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 109328 480 109356 2926
rect 110524 480 110552 2926
rect 111628 480 111656 4694
rect 112824 480 112852 6886
rect 113284 5302 113312 84166
rect 114572 5370 114600 84166
rect 115216 9042 115244 85478
rect 116044 78062 116072 87790
rect 116308 87774 116348 87802
rect 118056 87802 118084 88049
rect 118976 87802 119004 88049
rect 119896 87938 119924 88049
rect 117216 87790 117268 87796
rect 116320 85542 116348 87774
rect 117976 87774 118084 87802
rect 118896 87774 119004 87802
rect 119264 87910 119924 87938
rect 116308 85536 116360 85542
rect 116308 85478 116360 85484
rect 117976 84194 118004 87774
rect 118896 87258 118924 87774
rect 117332 84166 118004 84194
rect 118712 87230 118924 87258
rect 116032 78056 116084 78062
rect 116032 77998 116084 78004
rect 117228 32428 117280 32434
rect 117228 32370 117280 32376
rect 115204 9036 115256 9042
rect 115204 8978 115256 8984
rect 114560 5364 114612 5370
rect 114560 5306 114612 5312
rect 113272 5296 113324 5302
rect 113272 5238 113324 5244
rect 115204 5092 115256 5098
rect 115204 5034 115256 5040
rect 114008 2916 114060 2922
rect 114008 2858 114060 2864
rect 114020 480 114048 2858
rect 115216 480 115244 5034
rect 117240 3738 117268 32370
rect 117332 17338 117360 84166
rect 117320 17332 117372 17338
rect 117320 17274 117372 17280
rect 118712 6186 118740 87230
rect 119264 84194 119292 87910
rect 120816 87802 120844 88049
rect 121736 87802 121764 88049
rect 122656 87802 122684 88049
rect 123576 87802 123604 88049
rect 124496 87802 124524 88049
rect 125324 87802 125352 88049
rect 126244 87802 126272 88049
rect 127164 87802 127192 88049
rect 128084 87802 128112 88049
rect 129004 87802 129032 88049
rect 129924 87802 129952 88049
rect 130844 87938 130872 88049
rect 120816 87774 120856 87802
rect 120828 85542 120856 87774
rect 121656 87774 121764 87802
rect 122576 87774 122684 87802
rect 123496 87774 123604 87802
rect 124416 87774 124524 87802
rect 125244 87774 125352 87802
rect 126164 87774 126272 87802
rect 126992 87774 127192 87802
rect 128004 87774 128112 87802
rect 128924 87774 129032 87802
rect 129752 87774 129952 87802
rect 130304 87910 130872 87938
rect 121656 87258 121684 87774
rect 121472 87230 121684 87258
rect 119344 85536 119396 85542
rect 119344 85478 119396 85484
rect 120816 85536 120868 85542
rect 120816 85478 120868 85484
rect 118804 84166 119292 84194
rect 118804 18698 118832 84166
rect 118792 18692 118844 18698
rect 118792 18634 118844 18640
rect 119356 14482 119384 85478
rect 121472 24138 121500 87230
rect 122576 84194 122604 87774
rect 123496 84194 123524 87774
rect 124416 87122 124444 87774
rect 121564 84166 122604 84194
rect 122852 84166 123524 84194
rect 124232 87094 124444 87122
rect 121564 73846 121592 84166
rect 121552 73840 121604 73846
rect 121552 73782 121604 73788
rect 122852 26994 122880 84166
rect 122840 26988 122892 26994
rect 122840 26930 122892 26936
rect 124128 26512 124180 26518
rect 124128 26454 124180 26460
rect 121460 24132 121512 24138
rect 121460 24074 121512 24080
rect 119344 14476 119396 14482
rect 119344 14418 119396 14424
rect 119896 14476 119948 14482
rect 119896 14418 119948 14424
rect 118700 6180 118752 6186
rect 118700 6122 118752 6128
rect 118792 5024 118844 5030
rect 118792 4966 118844 4972
rect 116400 3732 116452 3738
rect 116400 3674 116452 3680
rect 117228 3732 117280 3738
rect 117228 3674 117280 3680
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 116412 480 116440 3674
rect 117608 480 117636 3674
rect 118804 480 118832 4966
rect 119908 480 119936 14418
rect 122288 4820 122340 4826
rect 122288 4762 122340 4768
rect 121092 2576 121144 2582
rect 121092 2518 121144 2524
rect 121104 480 121132 2518
rect 122300 480 122328 4762
rect 124140 3534 124168 26454
rect 124232 6254 124260 87094
rect 125244 84194 125272 87774
rect 126164 84194 126192 87774
rect 124324 84166 125272 84194
rect 125612 84166 126192 84194
rect 124324 8974 124352 84166
rect 125612 11830 125640 84166
rect 126992 21486 127020 87774
rect 128004 84194 128032 87774
rect 128924 84194 128952 87774
rect 127084 84166 128032 84194
rect 128372 84166 128952 84194
rect 127084 29646 127112 84166
rect 128372 32434 128400 84166
rect 129648 83496 129700 83502
rect 129648 83438 129700 83444
rect 128360 32428 128412 32434
rect 128360 32370 128412 32376
rect 127072 29640 127124 29646
rect 127072 29582 127124 29588
rect 128268 24268 128320 24274
rect 128268 24210 128320 24216
rect 126980 21480 127032 21486
rect 126980 21422 127032 21428
rect 125600 11824 125652 11830
rect 125600 11766 125652 11772
rect 128176 10464 128228 10470
rect 128176 10406 128228 10412
rect 124312 8968 124364 8974
rect 124312 8910 124364 8916
rect 124220 6248 124272 6254
rect 124220 6190 124272 6196
rect 125876 6180 125928 6186
rect 125876 6122 125928 6128
rect 124680 3732 124732 3738
rect 124680 3674 124732 3680
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 123496 480 123524 3470
rect 124692 480 124720 3674
rect 125888 480 125916 6122
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 10406
rect 128280 3534 128308 24210
rect 128268 3528 128320 3534
rect 128268 3470 128320 3476
rect 128360 2848 128412 2854
rect 128358 2816 128360 2825
rect 128412 2816 128414 2825
rect 129660 2774 129688 83438
rect 129752 14482 129780 87774
rect 130304 84194 130332 87910
rect 131764 87802 131792 88049
rect 132592 87802 132620 88049
rect 133512 87802 133540 88049
rect 134432 87802 134460 88049
rect 135352 87802 135380 88049
rect 136272 87802 136300 88049
rect 137192 87802 137220 88049
rect 138112 87802 138140 88049
rect 139032 87802 139060 88049
rect 139860 87802 139888 88049
rect 131764 87774 131804 87802
rect 132592 87774 132632 87802
rect 131776 85542 131804 87774
rect 130384 85536 130436 85542
rect 130384 85478 130436 85484
rect 131764 85536 131816 85542
rect 131764 85478 131816 85484
rect 129844 84166 130332 84194
rect 129844 26518 129872 84166
rect 130396 57254 130424 85478
rect 132604 85134 132632 87774
rect 133432 87774 133540 87802
rect 134352 87774 134460 87802
rect 135272 87774 135380 87802
rect 136192 87774 136300 87802
rect 137112 87774 137220 87802
rect 138032 87774 138140 87802
rect 138952 87774 139060 87802
rect 139780 87774 139888 87802
rect 140780 87802 140808 88049
rect 141700 87802 141728 88049
rect 142620 87802 142648 88049
rect 140780 87774 140912 87802
rect 141700 87774 141740 87802
rect 132592 85128 132644 85134
rect 132592 85070 132644 85076
rect 133432 84194 133460 87774
rect 134352 84194 134380 87774
rect 132604 84166 133460 84194
rect 133984 84166 134380 84194
rect 130384 57248 130436 57254
rect 130384 57190 130436 57196
rect 129832 26512 129884 26518
rect 129832 26454 129884 26460
rect 129740 14476 129792 14482
rect 129740 14418 129792 14424
rect 131764 11756 131816 11762
rect 131764 11698 131816 11704
rect 130568 8968 130620 8974
rect 130568 8910 130620 8916
rect 128358 2751 128414 2760
rect 129384 2746 129688 2774
rect 129384 480 129412 2746
rect 130580 480 130608 8910
rect 131776 480 131804 11698
rect 132222 2952 132278 2961
rect 132222 2887 132278 2896
rect 132236 2854 132264 2887
rect 132224 2848 132276 2854
rect 132604 2825 132632 84166
rect 133788 80776 133840 80782
rect 133788 80718 133840 80724
rect 133800 4078 133828 80718
rect 132960 4072 133012 4078
rect 132960 4014 133012 4020
rect 133788 4072 133840 4078
rect 133788 4014 133840 4020
rect 132224 2790 132276 2796
rect 132590 2816 132646 2825
rect 132590 2751 132646 2760
rect 132972 480 133000 4014
rect 133984 3602 134012 84166
rect 135168 35216 135220 35222
rect 135168 35158 135220 35164
rect 135180 4078 135208 35158
rect 134156 4072 134208 4078
rect 134156 4014 134208 4020
rect 135168 4072 135220 4078
rect 135168 4014 135220 4020
rect 133972 3596 134024 3602
rect 133972 3538 134024 3544
rect 134064 3596 134116 3602
rect 134064 3538 134116 3544
rect 134076 2961 134104 3538
rect 134062 2952 134118 2961
rect 134062 2887 134118 2896
rect 134168 480 134196 4014
rect 135272 3466 135300 87774
rect 136192 84194 136220 87774
rect 137112 84194 137140 87774
rect 135364 84166 136220 84194
rect 136652 84166 137140 84194
rect 135364 4214 135392 84166
rect 136548 14476 136600 14482
rect 136548 14418 136600 14424
rect 135444 11824 135496 11830
rect 135444 11766 135496 11772
rect 135352 4208 135404 4214
rect 135352 4150 135404 4156
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135456 2774 135484 11766
rect 136560 2774 136588 14418
rect 136652 3670 136680 84166
rect 137928 78056 137980 78062
rect 137928 77998 137980 78004
rect 136640 3664 136692 3670
rect 136640 3606 136692 3612
rect 137940 2774 137968 77998
rect 138032 3942 138060 87774
rect 138952 84194 138980 87774
rect 139780 84194 139808 87774
rect 140780 86148 140832 86154
rect 140780 86090 140832 86096
rect 138124 84166 138980 84194
rect 139412 84166 139808 84194
rect 138124 4010 138152 84166
rect 139308 14612 139360 14618
rect 139308 14554 139360 14560
rect 138112 4004 138164 4010
rect 138112 3946 138164 3952
rect 138020 3936 138072 3942
rect 138020 3878 138072 3884
rect 139320 3534 139348 14554
rect 139412 3602 139440 84166
rect 140792 42090 140820 86090
rect 140884 55894 140912 87774
rect 141712 86154 141740 87774
rect 142540 87774 142648 87802
rect 143540 87802 143568 88049
rect 144460 87802 144488 88049
rect 145380 87802 145408 88049
rect 143540 87774 143580 87802
rect 141700 86148 141752 86154
rect 141700 86090 141752 86096
rect 142540 84194 142568 87774
rect 142172 84166 142568 84194
rect 140872 55888 140924 55894
rect 140872 55830 140924 55836
rect 142172 53106 142200 84166
rect 143448 80708 143500 80714
rect 143448 80650 143500 80656
rect 142160 53100 142212 53106
rect 142160 53042 142212 53048
rect 140780 42084 140832 42090
rect 140780 42026 140832 42032
rect 142068 21412 142120 21418
rect 142068 21354 142120 21360
rect 140688 18692 140740 18698
rect 140688 18634 140740 18640
rect 139400 3596 139452 3602
rect 139400 3538 139452 3544
rect 140700 3534 140728 18634
rect 142080 3534 142108 21354
rect 143460 3534 143488 80650
rect 143552 47598 143580 87774
rect 144380 87774 144488 87802
rect 145300 87774 145408 87802
rect 146300 87802 146328 88049
rect 147128 87938 147156 88049
rect 146864 87910 147156 87938
rect 146300 87774 146340 87802
rect 144380 84194 144408 87774
rect 145300 84194 145328 87774
rect 143644 84166 144408 84194
rect 144932 84166 145328 84194
rect 143644 50386 143672 84166
rect 143632 50380 143684 50386
rect 143632 50322 143684 50328
rect 143540 47592 143592 47598
rect 143540 47534 143592 47540
rect 144932 44878 144960 84166
rect 146208 61396 146260 61402
rect 146208 61338 146260 61344
rect 144920 44872 144972 44878
rect 144920 44814 144972 44820
rect 144828 29708 144880 29714
rect 144828 29650 144880 29656
rect 144736 17332 144788 17338
rect 144736 17274 144788 17280
rect 144748 3602 144776 17274
rect 143540 3596 143592 3602
rect 143540 3538 143592 3544
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 135272 2746 135484 2774
rect 136468 2746 136588 2774
rect 137664 2746 137968 2774
rect 135272 480 135300 2746
rect 136468 480 136496 2746
rect 137664 480 137692 2746
rect 138860 480 138888 3470
rect 140056 480 140084 3470
rect 141252 480 141280 3470
rect 142448 480 142476 3470
rect 143552 480 143580 3538
rect 144840 3482 144868 29650
rect 146220 6914 146248 61338
rect 146312 39370 146340 87774
rect 146864 84194 146892 87910
rect 147772 87848 147824 87854
rect 147772 87790 147824 87796
rect 148048 87802 148076 88049
rect 148968 87854 148996 88049
rect 148956 87848 149008 87854
rect 146944 85536 146996 85542
rect 146944 85478 146996 85484
rect 146404 84166 146892 84194
rect 146404 75206 146432 84166
rect 146392 75200 146444 75206
rect 146392 75142 146444 75148
rect 146300 39364 146352 39370
rect 146300 39306 146352 39312
rect 146956 17270 146984 85478
rect 147588 21480 147640 21486
rect 147588 21422 147640 21428
rect 146944 17264 146996 17270
rect 146944 17206 146996 17212
rect 144748 3454 144868 3482
rect 145944 6886 146248 6914
rect 144748 480 144776 3454
rect 145944 480 145972 6886
rect 147600 3534 147628 21422
rect 147784 18630 147812 87790
rect 148048 87774 148088 87802
rect 149888 87802 149916 88049
rect 148956 87790 149008 87796
rect 148060 85542 148088 87774
rect 149808 87774 149916 87802
rect 150532 87848 150584 87854
rect 150808 87802 150836 88049
rect 151728 87854 151756 88049
rect 150532 87790 150584 87796
rect 148048 85536 148100 85542
rect 148048 85478 148100 85484
rect 149808 84194 149836 87774
rect 149072 84166 149836 84194
rect 148968 73908 149020 73914
rect 148968 73850 149020 73856
rect 147772 18624 147824 18630
rect 147772 18566 147824 18572
rect 148980 3534 149008 73850
rect 149072 4146 149100 84166
rect 150544 6914 150572 87790
rect 150728 87774 150836 87802
rect 151716 87848 151768 87854
rect 151716 87790 151768 87796
rect 152648 87802 152676 88049
rect 153568 87802 153596 88049
rect 154396 87802 154424 88049
rect 152648 87774 152688 87802
rect 150728 84194 150756 87774
rect 152660 85202 152688 87774
rect 153488 87774 153596 87802
rect 154316 87774 154424 87802
rect 155316 87802 155344 88049
rect 156236 87802 156264 88049
rect 157156 87802 157184 88049
rect 158076 87802 158104 88049
rect 155316 87774 155356 87802
rect 153488 86954 153516 87774
rect 153212 86926 153516 86954
rect 152648 85196 152700 85202
rect 152648 85138 152700 85144
rect 151728 85128 151780 85134
rect 151728 85070 151780 85076
rect 150452 6886 150572 6914
rect 150636 84166 150756 84194
rect 149060 4140 149112 4146
rect 149060 4082 149112 4088
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149520 3460 149572 3466
rect 149520 3402 149572 3408
rect 149532 480 149560 3402
rect 150452 3194 150480 6886
rect 150636 3618 150664 84166
rect 150544 3590 150664 3618
rect 150544 3398 150572 3590
rect 151740 3534 151768 85070
rect 153108 83564 153160 83570
rect 153108 83506 153160 83512
rect 153120 3534 153148 83506
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 150532 3392 150584 3398
rect 150532 3334 150584 3340
rect 150440 3188 150492 3194
rect 150440 3130 150492 3136
rect 150636 480 150664 3470
rect 151832 480 151860 3470
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 153212 3126 153240 86926
rect 154316 84194 154344 87774
rect 155328 85270 155356 87774
rect 156156 87774 156264 87802
rect 157076 87774 157184 87802
rect 157996 87774 158104 87802
rect 158720 87848 158772 87854
rect 158996 87802 159024 88049
rect 159916 87854 159944 88049
rect 158720 87790 158772 87796
rect 156156 86954 156184 87774
rect 155972 86926 156184 86954
rect 155316 85264 155368 85270
rect 155316 85206 155368 85212
rect 153304 84166 154344 84194
rect 153200 3120 153252 3126
rect 153200 3062 153252 3068
rect 153304 3058 153332 84166
rect 155868 75268 155920 75274
rect 155868 75210 155920 75216
rect 154212 3936 154264 3942
rect 154212 3878 154264 3884
rect 153292 3052 153344 3058
rect 153292 2994 153344 3000
rect 154224 480 154252 3878
rect 155880 3534 155908 75210
rect 155408 3528 155460 3534
rect 155408 3470 155460 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 155420 480 155448 3470
rect 155972 2990 156000 86926
rect 157076 84194 157104 87774
rect 157996 84194 158024 87774
rect 156064 84166 157104 84194
rect 157352 84166 158024 84194
rect 155960 2984 156012 2990
rect 155960 2926 156012 2932
rect 156064 2922 156092 84166
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 156052 2916 156104 2922
rect 156052 2858 156104 2864
rect 156616 480 156644 3538
rect 157352 2854 157380 84166
rect 157800 4004 157852 4010
rect 157800 3946 157852 3952
rect 157340 2848 157392 2854
rect 157340 2790 157392 2796
rect 157812 480 157840 3946
rect 158732 3738 158760 87790
rect 158916 87774 159024 87802
rect 159904 87848 159956 87854
rect 160836 87802 160864 88049
rect 159904 87790 159956 87796
rect 160756 87774 160864 87802
rect 161664 87802 161692 88049
rect 162584 87802 162612 88049
rect 163504 87802 163532 88049
rect 164424 87802 164452 88049
rect 161664 87774 161704 87802
rect 158916 84194 158944 87774
rect 160756 84194 160784 87774
rect 161388 85196 161440 85202
rect 161388 85138 161440 85144
rect 158824 84166 158944 84194
rect 160296 84166 160784 84194
rect 158720 3732 158772 3738
rect 158720 3674 158772 3680
rect 158824 3670 158852 84166
rect 160008 18760 160060 18766
rect 160008 18702 160060 18708
rect 160020 4146 160048 18702
rect 158904 4140 158956 4146
rect 158904 4082 158956 4088
rect 160008 4140 160060 4146
rect 160008 4082 160060 4088
rect 158812 3664 158864 3670
rect 158812 3606 158864 3612
rect 158916 480 158944 4082
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 160112 480 160140 3606
rect 160296 3505 160324 84166
rect 160282 3496 160338 3505
rect 160282 3431 160338 3440
rect 161400 2774 161428 85138
rect 161676 85066 161704 87774
rect 162504 87774 162612 87802
rect 163424 87774 163532 87802
rect 164344 87774 164452 87802
rect 165344 87802 165372 88049
rect 166264 87802 166292 88049
rect 165344 87774 165384 87802
rect 161664 85060 161716 85066
rect 161664 85002 161716 85008
rect 162504 84194 162532 87774
rect 163424 84194 163452 87774
rect 161584 84166 162532 84194
rect 162872 84166 163452 84194
rect 161584 3641 161612 84166
rect 162768 26988 162820 26994
rect 162768 26930 162820 26936
rect 161570 3632 161626 3641
rect 161570 3567 161626 3576
rect 162780 2774 162808 26930
rect 162872 3777 162900 84166
rect 163688 10532 163740 10538
rect 163688 10474 163740 10480
rect 162858 3768 162914 3777
rect 162858 3703 162914 3712
rect 161308 2746 161428 2774
rect 162504 2746 162808 2774
rect 161308 480 161336 2746
rect 162504 480 162532 2746
rect 163700 480 163728 10474
rect 164344 3369 164372 87774
rect 165356 84998 165384 87774
rect 166184 87774 166292 87802
rect 167000 87848 167052 87854
rect 167184 87802 167212 88049
rect 168104 87854 168132 88049
rect 167000 87790 167052 87796
rect 165344 84992 165396 84998
rect 165344 84934 165396 84940
rect 165528 84992 165580 84998
rect 165528 84934 165580 84940
rect 165540 4146 165568 84934
rect 166184 84194 166212 87774
rect 165632 84166 166212 84194
rect 165632 6186 165660 84166
rect 167012 80782 167040 87790
rect 167104 87774 167212 87802
rect 168092 87848 168144 87854
rect 168932 87802 168960 88049
rect 168092 87790 168144 87796
rect 168852 87774 168960 87802
rect 169760 87848 169812 87854
rect 169760 87790 169812 87796
rect 169852 87802 169880 88049
rect 170772 87854 170800 88049
rect 170760 87848 170812 87854
rect 167104 83502 167132 87774
rect 168852 84194 168880 87774
rect 168392 84166 168880 84194
rect 169024 84244 169076 84250
rect 169024 84186 169076 84192
rect 167092 83496 167144 83502
rect 167092 83438 167144 83444
rect 167000 80776 167052 80782
rect 167000 80718 167052 80724
rect 168392 14482 168420 84166
rect 169036 21486 169064 84186
rect 169024 21480 169076 21486
rect 169024 21422 169076 21428
rect 169772 17338 169800 87790
rect 169852 87774 169892 87802
rect 170760 87790 170812 87796
rect 171692 87802 171720 88049
rect 172612 87802 172640 88049
rect 173532 87802 173560 88049
rect 174452 87802 174480 88049
rect 171692 87774 171732 87802
rect 172612 87774 172652 87802
rect 169864 18698 169892 87774
rect 171704 84250 171732 87774
rect 172624 85134 172652 87774
rect 173452 87774 173560 87802
rect 174372 87774 174480 87802
rect 175372 87802 175400 88049
rect 176292 87802 176320 88049
rect 177120 87802 177148 88049
rect 178040 87802 178068 88049
rect 178960 87802 178988 88049
rect 179880 87802 179908 88049
rect 175372 87774 175412 87802
rect 176292 87774 176332 87802
rect 177120 87774 177160 87802
rect 178040 87774 178080 87802
rect 172612 85128 172664 85134
rect 172612 85070 172664 85076
rect 171692 84244 171744 84250
rect 173452 84194 173480 87774
rect 174372 84194 174400 87774
rect 175384 85202 175412 87774
rect 176016 85536 176068 85542
rect 176016 85478 176068 85484
rect 175924 85332 175976 85338
rect 175924 85274 175976 85280
rect 175372 85196 175424 85202
rect 175372 85138 175424 85144
rect 171692 84186 171744 84192
rect 172624 84166 173480 84194
rect 173912 84166 174400 84194
rect 169852 18692 169904 18698
rect 169852 18634 169904 18640
rect 169760 17332 169812 17338
rect 169760 17274 169812 17280
rect 168380 14476 168432 14482
rect 168380 14418 168432 14424
rect 170772 10668 170824 10674
rect 170772 10610 170824 10616
rect 168288 10600 168340 10606
rect 168288 10542 168340 10548
rect 166080 9036 166132 9042
rect 166080 8978 166132 8984
rect 165620 6180 165672 6186
rect 165620 6122 165672 6128
rect 164884 4140 164936 4146
rect 164884 4082 164936 4088
rect 165528 4140 165580 4146
rect 165528 4082 165580 4088
rect 164330 3360 164386 3369
rect 164330 3295 164386 3304
rect 164896 480 164924 4082
rect 166092 480 166120 8978
rect 168300 3398 168328 10542
rect 169576 9104 169628 9110
rect 169576 9046 169628 9052
rect 168380 3732 168432 3738
rect 168380 3674 168432 3680
rect 167184 3392 167236 3398
rect 167184 3334 167236 3340
rect 168288 3392 168340 3398
rect 168288 3334 168340 3340
rect 167196 480 167224 3334
rect 168392 480 168420 3674
rect 169588 480 169616 9046
rect 170784 480 170812 10610
rect 172624 3942 172652 84166
rect 173164 9172 173216 9178
rect 173164 9114 173216 9120
rect 172612 3936 172664 3942
rect 172612 3878 172664 3884
rect 171968 3188 172020 3194
rect 171968 3130 172020 3136
rect 171980 480 172008 3130
rect 173176 480 173204 9114
rect 173912 4010 173940 84166
rect 175188 10736 175240 10742
rect 175188 10678 175240 10684
rect 173900 4004 173952 4010
rect 173900 3946 173952 3952
rect 175200 3398 175228 10678
rect 174268 3392 174320 3398
rect 174268 3334 174320 3340
rect 175188 3392 175240 3398
rect 175188 3334 175240 3340
rect 175464 3392 175516 3398
rect 175464 3334 175516 3340
rect 174280 480 174308 3334
rect 175476 480 175504 3334
rect 175936 3194 175964 85274
rect 176028 3738 176056 85478
rect 176304 84998 176332 87774
rect 177132 85542 177160 87774
rect 177120 85536 177172 85542
rect 177120 85478 177172 85484
rect 178052 85338 178080 87774
rect 178880 87774 178988 87802
rect 179800 87774 179908 87802
rect 180800 87802 180828 88049
rect 181720 87802 181748 88049
rect 182640 87802 182668 88049
rect 183560 87802 183588 88049
rect 184388 87802 184416 88049
rect 185308 87802 185336 88049
rect 186228 87802 186256 88049
rect 180800 87774 180840 87802
rect 181720 87774 181760 87802
rect 182640 87774 182680 87802
rect 183560 87774 183600 87802
rect 184388 87774 184428 87802
rect 178040 85332 178092 85338
rect 178040 85274 178092 85280
rect 176292 84992 176344 84998
rect 176292 84934 176344 84940
rect 178880 84194 178908 87774
rect 179800 84194 179828 87774
rect 180812 85542 180840 87774
rect 180800 85536 180852 85542
rect 180800 85478 180852 85484
rect 178144 84166 178908 84194
rect 179432 84166 179828 84194
rect 181732 84194 181760 87774
rect 182652 85542 182680 87774
rect 182180 85536 182232 85542
rect 182180 85478 182232 85484
rect 182640 85536 182692 85542
rect 182640 85478 182692 85484
rect 181732 84166 182128 84194
rect 177856 10804 177908 10810
rect 177856 10746 177908 10752
rect 176660 9376 176712 9382
rect 176660 9318 176712 9324
rect 176016 3732 176068 3738
rect 176016 3674 176068 3680
rect 175924 3188 175976 3194
rect 175924 3130 175976 3136
rect 176672 480 176700 9318
rect 177868 480 177896 10746
rect 178144 3398 178172 84166
rect 179432 3482 179460 84166
rect 181996 11008 182048 11014
rect 181996 10950 182048 10956
rect 180248 9444 180300 9450
rect 180248 9386 180300 9392
rect 179064 3454 179460 3482
rect 178132 3392 178184 3398
rect 178132 3334 178184 3340
rect 179064 480 179092 3454
rect 180260 480 180288 9386
rect 182008 3398 182036 10950
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181996 3392 182048 3398
rect 181996 3334 182048 3340
rect 181456 480 181484 3334
rect 182100 3194 182128 84166
rect 182192 16574 182220 85478
rect 183572 85338 183600 87774
rect 184400 85542 184428 87774
rect 185228 87774 185336 87802
rect 186148 87774 186256 87802
rect 187148 87802 187176 88049
rect 188068 87802 188096 88049
rect 188988 87802 189016 88049
rect 187148 87774 187188 87802
rect 188068 87774 188108 87802
rect 184204 85536 184256 85542
rect 184204 85478 184256 85484
rect 184388 85536 184440 85542
rect 184388 85478 184440 85484
rect 183560 85332 183612 85338
rect 183560 85274 183612 85280
rect 182192 16546 182588 16574
rect 182088 3188 182140 3194
rect 182088 3130 182140 3136
rect 182560 480 182588 16546
rect 183744 9512 183796 9518
rect 183744 9454 183796 9460
rect 183756 480 183784 9454
rect 184216 5574 184244 85478
rect 184848 85332 184900 85338
rect 184848 85274 184900 85280
rect 184860 6322 184888 85274
rect 185228 84194 185256 87774
rect 186148 84194 186176 87774
rect 187160 85542 187188 87774
rect 188080 85542 188108 87774
rect 188908 87774 189016 87802
rect 189908 87802 189936 88049
rect 190828 87802 190856 88049
rect 191656 87802 191684 88049
rect 192576 87802 192604 88049
rect 193496 87802 193524 88049
rect 194416 87802 194444 88049
rect 195336 87802 195364 88049
rect 196256 87802 196284 88049
rect 197176 87802 197204 88049
rect 198096 87802 198124 88049
rect 198924 87802 198952 88049
rect 199844 87802 199872 88049
rect 200764 87802 200792 88049
rect 201684 87802 201712 88049
rect 202604 87802 202632 88049
rect 203524 87802 203552 88049
rect 204444 87802 204472 88049
rect 205364 87802 205392 88049
rect 206192 87802 206220 88049
rect 207112 87802 207140 88049
rect 208032 87802 208060 88049
rect 208952 87802 208980 88049
rect 209872 87802 209900 88049
rect 210792 87802 210820 88049
rect 211712 87802 211740 88049
rect 212632 87802 212660 88049
rect 213460 87802 213488 88049
rect 214380 87802 214408 88049
rect 215300 87802 215328 88049
rect 216220 87802 216248 88049
rect 217140 87802 217168 88049
rect 218060 87802 218088 88049
rect 218980 87802 219008 88049
rect 219900 87802 219928 88049
rect 220728 87802 220756 88049
rect 189908 87774 189948 87802
rect 190828 87774 190868 87802
rect 191656 87774 191788 87802
rect 192576 87774 192616 87802
rect 193496 87774 193536 87802
rect 194416 87774 194456 87802
rect 195336 87774 195376 87802
rect 196256 87774 196296 87802
rect 197176 87774 197308 87802
rect 198096 87774 198136 87802
rect 198924 87774 198964 87802
rect 199844 87774 199884 87802
rect 200764 87774 200804 87802
rect 201684 87774 201724 87802
rect 202604 87774 202644 87802
rect 203524 87774 203564 87802
rect 204444 87774 204484 87802
rect 205364 87774 205404 87802
rect 206192 87774 206232 87802
rect 207112 87774 207152 87802
rect 208032 87774 208072 87802
rect 208952 87774 208992 87802
rect 209872 87774 209912 87802
rect 210792 87774 210832 87802
rect 211712 87774 211752 87802
rect 212632 87774 212672 87802
rect 213460 87774 213500 87802
rect 214380 87774 214420 87802
rect 215300 87774 215340 87802
rect 216220 87774 216260 87802
rect 217140 87774 217180 87802
rect 218060 87774 218100 87802
rect 218980 87774 219020 87802
rect 219900 87774 219940 87802
rect 186964 85536 187016 85542
rect 186964 85478 187016 85484
rect 187148 85536 187200 85542
rect 187148 85478 187200 85484
rect 187608 85536 187660 85542
rect 187608 85478 187660 85484
rect 188068 85536 188120 85542
rect 188068 85478 188120 85484
rect 184952 84166 185256 84194
rect 186056 84166 186176 84194
rect 184952 83502 184980 84166
rect 184940 83496 184992 83502
rect 184940 83438 184992 83444
rect 184848 6316 184900 6322
rect 184848 6258 184900 6264
rect 184204 5568 184256 5574
rect 184204 5510 184256 5516
rect 186056 3942 186084 84166
rect 186976 14550 187004 85478
rect 186964 14544 187016 14550
rect 186964 14486 187016 14492
rect 186136 11892 186188 11898
rect 186136 11834 186188 11840
rect 186044 3936 186096 3942
rect 186044 3878 186096 3884
rect 186148 3398 186176 11834
rect 187332 9580 187384 9586
rect 187332 9522 187384 9528
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 186136 3392 186188 3398
rect 186136 3334 186188 3340
rect 184952 480 184980 3334
rect 186136 3188 186188 3194
rect 186136 3130 186188 3136
rect 186148 480 186176 3130
rect 187344 480 187372 9522
rect 187620 3738 187648 85478
rect 188908 18630 188936 87774
rect 188988 85536 189040 85542
rect 188988 85478 189040 85484
rect 188896 18624 188948 18630
rect 188896 18566 188948 18572
rect 188528 12096 188580 12102
rect 188528 12038 188580 12044
rect 187608 3732 187660 3738
rect 187608 3674 187660 3680
rect 188540 480 188568 12038
rect 189000 6254 189028 85478
rect 189920 84998 189948 87774
rect 190840 85542 190868 87774
rect 190828 85536 190880 85542
rect 190828 85478 190880 85484
rect 191656 85536 191708 85542
rect 191656 85478 191708 85484
rect 189908 84992 189960 84998
rect 189908 84934 189960 84940
rect 190828 9648 190880 9654
rect 190828 9590 190880 9596
rect 188988 6248 189040 6254
rect 188988 6190 189040 6196
rect 189724 5568 189776 5574
rect 189724 5510 189776 5516
rect 189736 480 189764 5510
rect 190840 480 190868 9590
rect 191668 6186 191696 85478
rect 191656 6180 191708 6186
rect 191656 6122 191708 6128
rect 191760 5166 191788 87774
rect 192588 85542 192616 87774
rect 193508 85542 193536 87774
rect 192576 85536 192628 85542
rect 192576 85478 192628 85484
rect 193128 85536 193180 85542
rect 193128 85478 193180 85484
rect 193496 85536 193548 85542
rect 193496 85478 193548 85484
rect 193036 12164 193088 12170
rect 193036 12106 193088 12112
rect 191748 5160 191800 5166
rect 191748 5102 191800 5108
rect 193048 2990 193076 12106
rect 193140 5098 193168 85478
rect 194428 16574 194456 87774
rect 195348 85542 195376 87774
rect 196268 85542 196296 87774
rect 194508 85536 194560 85542
rect 194508 85478 194560 85484
rect 195336 85536 195388 85542
rect 195336 85478 195388 85484
rect 195888 85536 195940 85542
rect 195888 85478 195940 85484
rect 196256 85536 196308 85542
rect 196256 85478 196308 85484
rect 197176 85536 197228 85542
rect 197176 85478 197228 85484
rect 194244 16546 194456 16574
rect 193220 6316 193272 6322
rect 193220 6258 193272 6264
rect 193128 5092 193180 5098
rect 193128 5034 193180 5040
rect 192024 2984 192076 2990
rect 192024 2926 192076 2932
rect 193036 2984 193088 2990
rect 193036 2926 193088 2932
rect 192036 480 192064 2926
rect 193232 480 193260 6258
rect 194244 4282 194272 16546
rect 194520 11778 194548 85478
rect 195244 84992 195296 84998
rect 195244 84934 195296 84940
rect 195256 14482 195284 84934
rect 195244 14476 195296 14482
rect 195244 14418 195296 14424
rect 195612 12232 195664 12238
rect 195612 12174 195664 12180
rect 194336 11750 194548 11778
rect 194232 4276 194284 4282
rect 194232 4218 194284 4224
rect 194336 4214 194364 11750
rect 194416 8900 194468 8906
rect 194416 8842 194468 8848
rect 194324 4208 194376 4214
rect 194324 4150 194376 4156
rect 194428 480 194456 8842
rect 195624 480 195652 12174
rect 195900 4486 195928 85478
rect 196808 14544 196860 14550
rect 196808 14486 196860 14492
rect 195888 4480 195940 4486
rect 195888 4422 195940 4428
rect 196820 480 196848 14486
rect 197188 4554 197216 85478
rect 197280 4622 197308 87774
rect 198108 85542 198136 87774
rect 198936 85542 198964 87774
rect 199856 87530 199884 87774
rect 199856 87502 200068 87530
rect 198096 85536 198148 85542
rect 198096 85478 198148 85484
rect 198648 85536 198700 85542
rect 198648 85478 198700 85484
rect 198924 85536 198976 85542
rect 198924 85478 198976 85484
rect 199936 85536 199988 85542
rect 199936 85478 199988 85484
rect 197912 8832 197964 8838
rect 197912 8774 197964 8780
rect 197268 4616 197320 4622
rect 197268 4558 197320 4564
rect 197176 4548 197228 4554
rect 197176 4490 197228 4496
rect 197924 480 197952 8774
rect 198660 4690 198688 85478
rect 199844 12300 199896 12306
rect 199844 12242 199896 12248
rect 198648 4684 198700 4690
rect 198648 4626 198700 4632
rect 199856 3194 199884 12242
rect 199948 4758 199976 85478
rect 200040 5370 200068 87502
rect 200776 85542 200804 87774
rect 201696 85542 201724 87774
rect 200764 85536 200816 85542
rect 200764 85478 200816 85484
rect 201408 85536 201460 85542
rect 201408 85478 201460 85484
rect 201684 85536 201736 85542
rect 201684 85478 201736 85484
rect 200120 83496 200172 83502
rect 200120 83438 200172 83444
rect 200132 16574 200160 83438
rect 200132 16546 200344 16574
rect 200028 5364 200080 5370
rect 200028 5306 200080 5312
rect 199936 4752 199988 4758
rect 199936 4694 199988 4700
rect 199108 3188 199160 3194
rect 199108 3130 199160 3136
rect 199844 3188 199896 3194
rect 199844 3130 199896 3136
rect 199120 480 199148 3130
rect 200316 480 200344 16546
rect 201420 5302 201448 85478
rect 202616 84194 202644 87774
rect 203536 85542 203564 87774
rect 204456 85542 204484 87774
rect 205376 86986 205404 87774
rect 205376 86958 205588 86986
rect 202788 85536 202840 85542
rect 202788 85478 202840 85484
rect 203524 85536 203576 85542
rect 203524 85478 203576 85484
rect 204168 85536 204220 85542
rect 204168 85478 204220 85484
rect 204444 85536 204496 85542
rect 204444 85478 204496 85484
rect 205456 85536 205508 85542
rect 205456 85478 205508 85484
rect 202616 84166 202736 84194
rect 202604 12368 202656 12374
rect 202604 12310 202656 12316
rect 201500 8628 201552 8634
rect 201500 8570 201552 8576
rect 201408 5296 201460 5302
rect 201408 5238 201460 5244
rect 201512 480 201540 8570
rect 202616 3482 202644 12310
rect 202708 4826 202736 84166
rect 202800 5234 202828 85478
rect 202788 5228 202840 5234
rect 202788 5170 202840 5176
rect 204180 5030 204208 85478
rect 205088 8560 205140 8566
rect 205088 8502 205140 8508
rect 204168 5024 204220 5030
rect 204168 4966 204220 4972
rect 202696 4820 202748 4826
rect 202696 4762 202748 4768
rect 203892 3936 203944 3942
rect 203892 3878 203944 3884
rect 202616 3454 202736 3482
rect 202708 480 202736 3454
rect 203904 480 203932 3878
rect 205100 480 205128 8502
rect 205272 5296 205324 5302
rect 205270 5264 205272 5273
rect 205324 5264 205326 5273
rect 205468 5234 205496 85478
rect 205560 5302 205588 86958
rect 206204 85542 206232 87774
rect 206192 85536 206244 85542
rect 206192 85478 206244 85484
rect 206928 85536 206980 85542
rect 206928 85478 206980 85484
rect 206940 32570 206968 85478
rect 207124 85338 207152 87774
rect 207112 85332 207164 85338
rect 207112 85274 207164 85280
rect 208044 84454 208072 87774
rect 208964 85542 208992 87774
rect 208952 85536 209004 85542
rect 208952 85478 209004 85484
rect 209688 85536 209740 85542
rect 209688 85478 209740 85484
rect 209044 85332 209096 85338
rect 209044 85274 209096 85280
rect 208032 84448 208084 84454
rect 208032 84390 208084 84396
rect 209056 35494 209084 85274
rect 209044 35488 209096 35494
rect 209044 35430 209096 35436
rect 206928 32564 206980 32570
rect 206928 32506 206980 32512
rect 209700 17338 209728 85478
rect 209884 85338 209912 87774
rect 209872 85332 209924 85338
rect 209872 85274 209924 85280
rect 210804 84194 210832 87774
rect 211724 85542 211752 87774
rect 212644 85542 212672 87774
rect 211712 85536 211764 85542
rect 211712 85478 211764 85484
rect 212448 85536 212500 85542
rect 212448 85478 212500 85484
rect 212632 85536 212684 85542
rect 212632 85478 212684 85484
rect 211804 84448 211856 84454
rect 211804 84390 211856 84396
rect 210804 84166 211108 84194
rect 211080 42158 211108 84166
rect 211068 42152 211120 42158
rect 211068 42094 211120 42100
rect 211816 38214 211844 84390
rect 212460 44946 212488 85478
rect 213472 84194 213500 87774
rect 214392 85542 214420 87774
rect 215312 85542 215340 87774
rect 213828 85536 213880 85542
rect 213828 85478 213880 85484
rect 214380 85536 214432 85542
rect 214380 85478 214432 85484
rect 215208 85536 215260 85542
rect 215208 85478 215260 85484
rect 215300 85536 215352 85542
rect 215300 85478 215352 85484
rect 213472 84166 213776 84194
rect 213748 50454 213776 84166
rect 213736 50448 213788 50454
rect 213736 50390 213788 50396
rect 213840 47666 213868 85478
rect 214564 85332 214616 85338
rect 214564 85274 214616 85280
rect 213828 47660 213880 47666
rect 213828 47602 213880 47608
rect 212448 44940 212500 44946
rect 212448 44882 212500 44888
rect 214576 39438 214604 85274
rect 215220 53242 215248 85478
rect 216232 84194 216260 87774
rect 217152 85542 217180 87774
rect 218072 85542 218100 87774
rect 216588 85536 216640 85542
rect 216588 85478 216640 85484
rect 217140 85536 217192 85542
rect 217140 85478 217192 85484
rect 217968 85536 218020 85542
rect 217968 85478 218020 85484
rect 218060 85536 218112 85542
rect 218060 85478 218112 85484
rect 216232 84166 216536 84194
rect 216508 57390 216536 84166
rect 216496 57384 216548 57390
rect 216496 57326 216548 57332
rect 216600 56166 216628 85478
rect 217980 60178 218008 85478
rect 218992 84194 219020 87774
rect 219912 85542 219940 87774
rect 220648 87774 220756 87802
rect 221648 87802 221676 88049
rect 222568 87802 222596 88049
rect 223488 87802 223516 88049
rect 221648 87774 221688 87802
rect 222568 87774 222608 87802
rect 219348 85536 219400 85542
rect 219348 85478 219400 85484
rect 219900 85536 219952 85542
rect 219900 85478 219952 85484
rect 218992 84166 219296 84194
rect 219268 65618 219296 84166
rect 219256 65612 219308 65618
rect 219256 65554 219308 65560
rect 219360 62966 219388 85478
rect 220648 71126 220676 87774
rect 220728 85536 220780 85542
rect 220728 85478 220780 85484
rect 220636 71120 220688 71126
rect 220636 71062 220688 71068
rect 220740 68406 220768 85478
rect 221660 85338 221688 87774
rect 222580 85542 222608 87774
rect 223408 87774 223516 87802
rect 224408 87802 224436 88049
rect 225328 87802 225356 88049
rect 226248 87802 226276 88049
rect 227168 87802 227196 88049
rect 227996 87802 228024 88049
rect 228916 87802 228944 88049
rect 229836 87802 229864 88049
rect 230756 87802 230784 88049
rect 231676 87802 231704 88049
rect 232596 87802 232624 88049
rect 233516 87802 233544 88049
rect 234436 87802 234464 88049
rect 235264 87802 235292 88049
rect 236184 87802 236212 88049
rect 237104 87938 237132 88049
rect 237104 87910 237328 87938
rect 224408 87774 224448 87802
rect 225328 87774 225368 87802
rect 226248 87774 226288 87802
rect 227168 87774 227208 87802
rect 227996 87774 228036 87802
rect 228916 87774 228956 87802
rect 229836 87774 229876 87802
rect 230756 87774 230796 87802
rect 231676 87774 231716 87802
rect 232596 87774 232636 87802
rect 233516 87774 233556 87802
rect 234436 87774 234568 87802
rect 235264 87774 235304 87802
rect 236184 87774 236224 87802
rect 222568 85536 222620 85542
rect 222568 85478 222620 85484
rect 221648 85332 221700 85338
rect 221648 85274 221700 85280
rect 220728 68400 220780 68406
rect 220728 68342 220780 68348
rect 219348 62960 219400 62966
rect 219348 62902 219400 62908
rect 217968 60172 218020 60178
rect 217968 60114 218020 60120
rect 216588 56160 216640 56166
rect 216588 56102 216640 56108
rect 215208 53236 215260 53242
rect 215208 53178 215260 53184
rect 214564 39432 214616 39438
rect 214564 39374 214616 39380
rect 211804 38208 211856 38214
rect 211804 38150 211856 38156
rect 223304 29776 223356 29782
rect 223304 29718 223356 29724
rect 213920 18624 213972 18630
rect 213920 18566 213972 18572
rect 209688 17332 209740 17338
rect 209688 17274 209740 17280
rect 213932 16574 213960 18566
rect 213932 16546 214512 16574
rect 206928 12436 206980 12442
rect 206928 12378 206980 12384
rect 205548 5296 205600 5302
rect 205548 5238 205600 5244
rect 205270 5199 205326 5208
rect 205364 5228 205416 5234
rect 205364 5170 205416 5176
rect 205456 5228 205508 5234
rect 205456 5170 205508 5176
rect 205376 5137 205404 5170
rect 205362 5128 205418 5137
rect 205362 5063 205418 5072
rect 206940 3398 206968 12378
rect 211068 11688 211120 11694
rect 211068 11630 211120 11636
rect 208584 8492 208636 8498
rect 208584 8434 208636 8440
rect 207388 3732 207440 3738
rect 207388 3674 207440 3680
rect 206192 3392 206244 3398
rect 206192 3334 206244 3340
rect 206928 3392 206980 3398
rect 206928 3334 206980 3340
rect 206204 480 206232 3334
rect 207400 480 207428 3674
rect 208596 480 208624 8434
rect 210976 6248 211028 6254
rect 210976 6190 211028 6196
rect 209686 5264 209742 5273
rect 209686 5199 209742 5208
rect 209594 5128 209650 5137
rect 209594 5063 209650 5072
rect 209608 4826 209636 5063
rect 209700 5030 209728 5199
rect 209688 5024 209740 5030
rect 209688 4966 209740 4972
rect 209596 4820 209648 4826
rect 209596 4762 209648 4768
rect 209780 3392 209832 3398
rect 209780 3334 209832 3340
rect 209792 480 209820 3334
rect 210988 480 211016 6190
rect 211080 3398 211108 11630
rect 213828 11620 213880 11626
rect 213828 11562 213880 11568
rect 212172 8424 212224 8430
rect 212172 8366 212224 8372
rect 211068 3392 211120 3398
rect 211068 3334 211120 3340
rect 212184 480 212212 8366
rect 213840 3398 213868 11562
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 213380 480 213408 3334
rect 214484 480 214512 16546
rect 218060 14476 218112 14482
rect 218060 14418 218112 14424
rect 217968 11552 218020 11558
rect 217968 11494 218020 11500
rect 215668 8356 215720 8362
rect 215668 8298 215720 8304
rect 215680 480 215708 8298
rect 217980 3398 218008 11494
rect 216864 3392 216916 3398
rect 216864 3334 216916 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 216876 480 216904 3334
rect 218072 480 218100 14418
rect 220452 11348 220504 11354
rect 220452 11290 220504 11296
rect 219256 8288 219308 8294
rect 219256 8230 219308 8236
rect 219268 480 219296 8230
rect 219440 5160 219492 5166
rect 219438 5128 219440 5137
rect 219492 5128 219494 5137
rect 219438 5063 219494 5072
rect 220464 480 220492 11290
rect 221556 6180 221608 6186
rect 221556 6122 221608 6128
rect 221568 480 221596 6122
rect 223316 3398 223344 29718
rect 223408 6458 223436 87774
rect 224420 85542 224448 87774
rect 225340 85542 225368 87774
rect 223488 85536 223540 85542
rect 223488 85478 223540 85484
rect 224408 85536 224460 85542
rect 224408 85478 224460 85484
rect 224868 85536 224920 85542
rect 224868 85478 224920 85484
rect 225328 85536 225380 85542
rect 225328 85478 225380 85484
rect 226156 85536 226208 85542
rect 226156 85478 226208 85484
rect 223500 6662 223528 85478
rect 224224 85332 224276 85338
rect 224224 85274 224276 85280
rect 224236 74118 224264 85274
rect 224224 74112 224276 74118
rect 224224 74054 224276 74060
rect 224776 11280 224828 11286
rect 224776 11222 224828 11228
rect 223488 6656 223540 6662
rect 223488 6598 223540 6604
rect 223396 6452 223448 6458
rect 223396 6394 223448 6400
rect 224788 3398 224816 11222
rect 224880 6390 224908 85478
rect 224868 6384 224920 6390
rect 224868 6326 224920 6332
rect 226168 6322 226196 85478
rect 226156 6316 226208 6322
rect 226156 6258 226208 6264
rect 226260 6254 226288 87774
rect 227180 85542 227208 87774
rect 227168 85536 227220 85542
rect 227168 85478 227220 85484
rect 227628 85536 227680 85542
rect 227628 85478 227680 85484
rect 227536 75336 227588 75342
rect 227536 75278 227588 75284
rect 227444 11212 227496 11218
rect 227444 11154 227496 11160
rect 226248 6248 226300 6254
rect 226248 6190 226300 6196
rect 225142 5128 225198 5137
rect 225142 5063 225198 5072
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 223304 3392 223356 3398
rect 223304 3334 223356 3340
rect 223948 3392 224000 3398
rect 223948 3334 224000 3340
rect 224776 3392 224828 3398
rect 224776 3334 224828 3340
rect 222764 480 222792 3334
rect 223960 480 223988 3334
rect 225156 480 225184 5063
rect 226340 3732 226392 3738
rect 226340 3674 226392 3680
rect 226352 480 226380 3674
rect 227456 3482 227484 11154
rect 227548 3738 227576 75278
rect 227640 6186 227668 85478
rect 228008 84658 228036 87774
rect 228928 84998 228956 87774
rect 229848 85542 229876 87774
rect 230768 85542 230796 87774
rect 229836 85536 229888 85542
rect 229836 85478 229888 85484
rect 230296 85536 230348 85542
rect 230296 85478 230348 85484
rect 230756 85536 230808 85542
rect 230756 85478 230808 85484
rect 228916 84992 228968 84998
rect 228916 84934 228968 84940
rect 227996 84652 228048 84658
rect 227996 84594 228048 84600
rect 229744 84652 229796 84658
rect 229744 84594 229796 84600
rect 229756 32502 229784 84594
rect 230308 39370 230336 85478
rect 230388 78124 230440 78130
rect 230388 78066 230440 78072
rect 230296 39364 230348 39370
rect 230296 39306 230348 39312
rect 229744 32496 229796 32502
rect 229744 32438 229796 32444
rect 227628 6180 227680 6186
rect 227628 6122 227680 6128
rect 228732 4140 228784 4146
rect 228732 4082 228784 4088
rect 227536 3732 227588 3738
rect 227536 3674 227588 3680
rect 227456 3454 227576 3482
rect 227548 480 227576 3454
rect 228744 480 228772 4082
rect 230400 3398 230428 78066
rect 231688 44878 231716 87774
rect 232608 85542 232636 87774
rect 233528 85542 233556 87774
rect 231768 85536 231820 85542
rect 231768 85478 231820 85484
rect 232596 85536 232648 85542
rect 232596 85478 232648 85484
rect 233148 85536 233200 85542
rect 233148 85478 233200 85484
rect 233516 85536 233568 85542
rect 233516 85478 233568 85484
rect 234436 85536 234488 85542
rect 234436 85478 234488 85484
rect 231676 44872 231728 44878
rect 231676 44814 231728 44820
rect 231676 43444 231728 43450
rect 231676 43386 231728 43392
rect 231688 3398 231716 43386
rect 231780 42090 231808 85478
rect 232504 84992 232556 84998
rect 232504 84934 232556 84940
rect 231768 42084 231820 42090
rect 231768 42026 231820 42032
rect 232516 38010 232544 84934
rect 233160 47598 233188 85478
rect 234448 50386 234476 85478
rect 234436 50380 234488 50386
rect 234436 50322 234488 50328
rect 233148 47592 233200 47598
rect 233148 47534 233200 47540
rect 232504 38004 232556 38010
rect 232504 37946 232556 37952
rect 234436 22976 234488 22982
rect 234436 22918 234488 22924
rect 232228 4208 232280 4214
rect 232228 4150 232280 4156
rect 229836 3392 229888 3398
rect 229836 3334 229888 3340
rect 230388 3392 230440 3398
rect 230388 3334 230440 3340
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231676 3392 231728 3398
rect 231676 3334 231728 3340
rect 229848 480 229876 3334
rect 231044 480 231072 3334
rect 232240 480 232268 4150
rect 234448 3398 234476 22918
rect 234540 14550 234568 87774
rect 235276 85542 235304 87774
rect 236196 85542 236224 87774
rect 235264 85536 235316 85542
rect 235264 85478 235316 85484
rect 235908 85536 235960 85542
rect 235908 85478 235960 85484
rect 236184 85536 236236 85542
rect 236184 85478 236236 85484
rect 237196 85536 237248 85542
rect 237196 85478 237248 85484
rect 235816 54528 235868 54534
rect 235816 54470 235868 54476
rect 234528 14544 234580 14550
rect 234528 14486 234580 14492
rect 235724 4276 235776 4282
rect 235724 4218 235776 4224
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 234436 3392 234488 3398
rect 234436 3334 234488 3340
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 233436 480 233464 3334
rect 234632 480 234660 3334
rect 235736 2122 235764 4218
rect 235828 3398 235856 54470
rect 235920 53106 235948 85478
rect 237208 55894 237236 85478
rect 237196 55888 237248 55894
rect 237196 55830 237248 55836
rect 235908 53100 235960 53106
rect 235908 53042 235960 53048
rect 237196 31136 237248 31142
rect 237196 31078 237248 31084
rect 237208 6914 237236 31078
rect 237300 18698 237328 87910
rect 238024 87802 238052 88049
rect 238944 87802 238972 88049
rect 239864 87802 239892 88049
rect 240784 87802 240812 88049
rect 241704 87802 241732 88049
rect 242532 87802 242560 88049
rect 243452 87802 243480 88049
rect 244372 87802 244400 88049
rect 245292 87802 245320 88049
rect 246212 87802 246240 88049
rect 247132 87802 247160 88049
rect 248052 87802 248080 88049
rect 248972 87802 249000 88049
rect 249800 87802 249828 88049
rect 250720 87802 250748 88049
rect 251640 87802 251668 88049
rect 252560 87802 252588 88049
rect 253480 87802 253508 88049
rect 254400 87802 254428 88049
rect 255320 87802 255348 88049
rect 256240 87802 256268 88049
rect 257068 87802 257096 88049
rect 257988 87802 258016 88049
rect 258908 87802 258936 88049
rect 259828 87802 259856 88049
rect 260748 87802 260776 88049
rect 238024 87774 238064 87802
rect 238944 87774 238984 87802
rect 239864 87774 239904 87802
rect 240784 87774 240824 87802
rect 241704 87774 241744 87802
rect 242532 87774 242572 87802
rect 243452 87774 243492 87802
rect 244372 87774 244412 87802
rect 245292 87774 245332 87802
rect 246212 87774 246252 87802
rect 247132 87774 247172 87802
rect 248052 87774 248092 87802
rect 248972 87774 249012 87802
rect 249800 87774 249840 87802
rect 250720 87774 250760 87802
rect 251640 87774 251680 87802
rect 252560 87774 252600 87802
rect 253480 87774 253520 87802
rect 254400 87774 254440 87802
rect 255320 87774 255360 87802
rect 256240 87774 256280 87802
rect 257068 87774 257108 87802
rect 257988 87774 258028 87802
rect 258908 87774 258948 87802
rect 259828 87774 259868 87802
rect 238036 85542 238064 87774
rect 238024 85536 238076 85542
rect 238024 85478 238076 85484
rect 238668 85536 238720 85542
rect 238668 85478 238720 85484
rect 238680 57254 238708 85478
rect 238956 85338 238984 87774
rect 238944 85332 238996 85338
rect 238944 85274 238996 85280
rect 239876 84998 239904 87774
rect 240796 85542 240824 87774
rect 241716 85542 241744 87774
rect 242544 87258 242572 87774
rect 242544 87230 242848 87258
rect 240784 85536 240836 85542
rect 240784 85478 240836 85484
rect 241336 85536 241388 85542
rect 241336 85478 241388 85484
rect 241704 85536 241756 85542
rect 241704 85478 241756 85484
rect 242716 85536 242768 85542
rect 242716 85478 242768 85484
rect 240784 85332 240836 85338
rect 240784 85274 240836 85280
rect 239864 84992 239916 84998
rect 239864 84934 239916 84940
rect 238668 57248 238720 57254
rect 238668 57190 238720 57196
rect 237288 18692 237340 18698
rect 237288 18634 237340 18640
rect 240796 13190 240824 85274
rect 241348 62830 241376 85478
rect 241428 80844 241480 80850
rect 241428 80786 241480 80792
rect 241336 62824 241388 62830
rect 241336 62766 241388 62772
rect 240784 13184 240836 13190
rect 240784 13126 240836 13132
rect 238668 11144 238720 11150
rect 238668 11086 238720 11092
rect 237024 6886 237236 6914
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 235736 2094 235856 2122
rect 235828 480 235856 2094
rect 237024 480 237052 6886
rect 238680 3398 238708 11086
rect 239312 4480 239364 4486
rect 239312 4422 239364 4428
rect 238116 3392 238168 3398
rect 238116 3334 238168 3340
rect 238668 3392 238720 3398
rect 238668 3334 238720 3340
rect 238128 480 238156 3334
rect 239324 480 239352 4422
rect 241440 3398 241468 80786
rect 242624 33856 242676 33862
rect 242624 33798 242676 33804
rect 242636 3398 242664 33798
rect 242728 21486 242756 85478
rect 242716 21480 242768 21486
rect 242716 21422 242768 21428
rect 242820 7478 242848 87230
rect 243464 85542 243492 87774
rect 244384 85542 244412 87774
rect 243452 85536 243504 85542
rect 243452 85478 243504 85484
rect 244188 85536 244240 85542
rect 244188 85478 244240 85484
rect 244372 85536 244424 85542
rect 244372 85478 244424 85484
rect 244096 25696 244148 25702
rect 244096 25638 244148 25644
rect 242808 7472 242860 7478
rect 242808 7414 242860 7420
rect 242900 4548 242952 4554
rect 242900 4490 242952 4496
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 241428 3392 241480 3398
rect 241428 3334 241480 3340
rect 241704 3392 241756 3398
rect 241704 3334 241756 3340
rect 242624 3392 242676 3398
rect 242624 3334 242676 3340
rect 240520 480 240548 3334
rect 241716 480 241744 3334
rect 242912 480 242940 4490
rect 244108 480 244136 25638
rect 244200 7546 244228 85478
rect 245304 84194 245332 87774
rect 246224 85542 246252 87774
rect 247144 85542 247172 87774
rect 245568 85536 245620 85542
rect 245568 85478 245620 85484
rect 246212 85536 246264 85542
rect 246212 85478 246264 85484
rect 246948 85536 247000 85542
rect 246948 85478 247000 85484
rect 247132 85536 247184 85542
rect 247132 85478 247184 85484
rect 245304 84166 245516 84194
rect 245384 36576 245436 36582
rect 245384 36518 245436 36524
rect 244188 7540 244240 7546
rect 244188 7482 244240 7488
rect 245396 6914 245424 36518
rect 245488 7750 245516 84166
rect 245580 8090 245608 85478
rect 245568 8084 245620 8090
rect 245568 8026 245620 8032
rect 246960 8022 246988 85478
rect 248064 84194 248092 87774
rect 248984 85542 249012 87774
rect 249812 85542 249840 87774
rect 248328 85536 248380 85542
rect 248328 85478 248380 85484
rect 248972 85536 249024 85542
rect 248972 85478 249024 85484
rect 249708 85536 249760 85542
rect 249708 85478 249760 85484
rect 249800 85536 249852 85542
rect 249800 85478 249852 85484
rect 248064 84166 248276 84194
rect 248144 28416 248196 28422
rect 248144 28358 248196 28364
rect 246948 8016 247000 8022
rect 246948 7958 247000 7964
rect 245476 7744 245528 7750
rect 245476 7686 245528 7692
rect 245212 6886 245424 6914
rect 245212 480 245240 6886
rect 246396 4616 246448 4622
rect 246396 4558 246448 4564
rect 246408 480 246436 4558
rect 248156 3398 248184 28358
rect 248248 7886 248276 84166
rect 248340 7954 248368 85478
rect 249064 84992 249116 84998
rect 249064 84934 249116 84940
rect 249076 60042 249104 84934
rect 249064 60036 249116 60042
rect 249064 59978 249116 59984
rect 249616 40724 249668 40730
rect 249616 40666 249668 40672
rect 248878 8936 248934 8945
rect 248878 8871 248934 8880
rect 248892 8294 248920 8871
rect 248880 8288 248932 8294
rect 248880 8230 248932 8236
rect 248328 7948 248380 7954
rect 248328 7890 248380 7896
rect 248236 7880 248288 7886
rect 248236 7822 248288 7828
rect 249628 3398 249656 40666
rect 249720 7410 249748 85478
rect 250732 84194 250760 87774
rect 251652 85542 251680 87774
rect 252572 85542 252600 87774
rect 251088 85536 251140 85542
rect 251088 85478 251140 85484
rect 251640 85536 251692 85542
rect 251640 85478 251692 85484
rect 252468 85536 252520 85542
rect 252468 85478 252520 85484
rect 252560 85536 252612 85542
rect 252560 85478 252612 85484
rect 250732 84166 251036 84194
rect 251008 15910 251036 84166
rect 250996 15904 251048 15910
rect 250996 15846 251048 15852
rect 251100 7818 251128 85478
rect 252284 67040 252336 67046
rect 252284 66982 252336 66988
rect 251088 7812 251140 7818
rect 251088 7754 251140 7760
rect 249708 7404 249760 7410
rect 249708 7346 249760 7352
rect 249984 4684 250036 4690
rect 249984 4626 250036 4632
rect 247592 3392 247644 3398
rect 247592 3334 247644 3340
rect 248144 3392 248196 3398
rect 248144 3334 248196 3340
rect 248788 3392 248840 3398
rect 248788 3334 248840 3340
rect 249616 3392 249668 3398
rect 249616 3334 249668 3340
rect 247604 480 247632 3334
rect 248800 480 248828 3334
rect 249996 480 250024 4626
rect 251180 3732 251232 3738
rect 251180 3674 251232 3680
rect 251192 480 251220 3674
rect 252296 3482 252324 66982
rect 252480 65550 252508 85478
rect 253492 84194 253520 87774
rect 254412 85542 254440 87774
rect 255332 85542 255360 87774
rect 253848 85536 253900 85542
rect 253848 85478 253900 85484
rect 254400 85536 254452 85542
rect 254400 85478 254452 85484
rect 255228 85536 255280 85542
rect 255228 85478 255280 85484
rect 255320 85536 255372 85542
rect 255320 85478 255372 85484
rect 253492 84166 253796 84194
rect 253768 68338 253796 84166
rect 253756 68332 253808 68338
rect 253756 68274 253808 68280
rect 252468 65544 252520 65550
rect 252468 65486 252520 65492
rect 253860 19990 253888 85478
rect 254584 84992 254636 84998
rect 254584 84934 254636 84940
rect 254596 21418 254624 84934
rect 255240 71058 255268 85478
rect 256252 84194 256280 87774
rect 256608 85536 256660 85542
rect 256608 85478 256660 85484
rect 256700 85536 256752 85542
rect 256700 85478 256752 85484
rect 256252 84166 256556 84194
rect 255228 71052 255280 71058
rect 255228 70994 255280 71000
rect 256424 46368 256476 46374
rect 256424 46310 256476 46316
rect 254584 21412 254636 21418
rect 254584 21354 254636 21360
rect 253848 19984 253900 19990
rect 253848 19926 253900 19932
rect 252376 10260 252428 10266
rect 252376 10202 252428 10208
rect 252388 3738 252416 10202
rect 255228 10192 255280 10198
rect 255228 10134 255280 10140
rect 253480 4752 253532 4758
rect 253480 4694 253532 4700
rect 252376 3732 252428 3738
rect 252376 3674 252428 3680
rect 252296 3454 252416 3482
rect 252388 480 252416 3454
rect 253492 480 253520 4694
rect 255240 3398 255268 10134
rect 256436 3398 256464 46310
rect 256528 37942 256556 84166
rect 256516 37936 256568 37942
rect 256516 37878 256568 37884
rect 256620 32434 256648 85478
rect 256712 83502 256740 85478
rect 257080 84250 257108 87774
rect 258000 85542 258028 87774
rect 258920 85542 258948 87774
rect 259840 85542 259868 87774
rect 260668 87774 260776 87802
rect 261668 87802 261696 88049
rect 262588 87802 262616 88049
rect 263508 87802 263536 88049
rect 261668 87774 261708 87802
rect 262588 87774 262628 87802
rect 257988 85536 258040 85542
rect 257988 85478 258040 85484
rect 258080 85536 258132 85542
rect 258080 85478 258132 85484
rect 258908 85536 258960 85542
rect 258908 85478 258960 85484
rect 259828 85536 259880 85542
rect 259828 85478 259880 85484
rect 257068 84244 257120 84250
rect 257068 84186 257120 84192
rect 256700 83496 256752 83502
rect 256700 83438 256752 83444
rect 258092 80782 258120 85478
rect 258724 84244 258776 84250
rect 258724 84186 258776 84192
rect 258080 80776 258132 80782
rect 258080 80718 258132 80724
rect 256608 32428 256660 32434
rect 256608 32370 256660 32376
rect 258736 14482 258764 84186
rect 260564 24200 260616 24206
rect 260564 24142 260616 24148
rect 258724 14476 258776 14482
rect 258724 14418 258776 14424
rect 259368 10124 259420 10130
rect 259368 10066 259420 10072
rect 257068 5364 257120 5370
rect 257068 5306 257120 5312
rect 254676 3392 254728 3398
rect 254676 3334 254728 3340
rect 255228 3392 255280 3398
rect 255228 3334 255280 3340
rect 255872 3392 255924 3398
rect 255872 3334 255924 3340
rect 256424 3392 256476 3398
rect 256424 3334 256476 3340
rect 254688 480 254716 3334
rect 255884 480 255912 3334
rect 257080 480 257108 5306
rect 259380 2990 259408 10066
rect 260576 3398 260604 24142
rect 260668 18630 260696 87774
rect 260748 85536 260800 85542
rect 260748 85478 260800 85484
rect 260656 18624 260708 18630
rect 260656 18566 260708 18572
rect 260760 17270 260788 85478
rect 261680 85338 261708 87774
rect 262600 85542 262628 87774
rect 263428 87774 263536 87802
rect 264336 87802 264364 88049
rect 265256 87802 265284 88049
rect 266176 87802 266204 88049
rect 267096 87802 267124 88049
rect 268016 87802 268044 88049
rect 268936 87802 268964 88049
rect 269856 87802 269884 88049
rect 270776 87802 270804 88049
rect 271604 87802 271632 88049
rect 272524 87802 272552 88049
rect 273444 87802 273472 88049
rect 274364 87802 274392 88049
rect 275284 87802 275312 88049
rect 276204 87802 276232 88049
rect 277124 87802 277152 88049
rect 278044 87802 278072 88049
rect 278964 87802 278992 88049
rect 279792 87802 279820 88049
rect 280712 87802 280740 88049
rect 281632 87802 281660 88049
rect 282552 87802 282580 88049
rect 283472 87802 283500 88049
rect 284392 87802 284420 88049
rect 285312 87802 285340 88049
rect 264336 87774 264376 87802
rect 265256 87774 265296 87802
rect 266176 87774 266216 87802
rect 267096 87774 267136 87802
rect 268016 87774 268056 87802
rect 268936 87774 268976 87802
rect 269856 87774 269896 87802
rect 270776 87774 270816 87802
rect 271604 87774 271644 87802
rect 272524 87774 272564 87802
rect 273444 87774 273484 87802
rect 274364 87774 274404 87802
rect 275284 87774 275324 87802
rect 276204 87774 276244 87802
rect 277124 87774 277164 87802
rect 278044 87774 278084 87802
rect 278964 87774 279004 87802
rect 279792 87774 279832 87802
rect 280712 87774 280752 87802
rect 281632 87774 281672 87802
rect 282552 87774 282592 87802
rect 262588 85536 262640 85542
rect 262588 85478 262640 85484
rect 261668 85332 261720 85338
rect 261668 85274 261720 85280
rect 263324 49088 263376 49094
rect 263324 49030 263376 49036
rect 260748 17264 260800 17270
rect 260748 17206 260800 17212
rect 261760 10056 261812 10062
rect 261760 9998 261812 10004
rect 260656 5024 260708 5030
rect 260656 4966 260708 4972
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 260564 3392 260616 3398
rect 260564 3334 260616 3340
rect 258264 2984 258316 2990
rect 258264 2926 258316 2932
rect 259368 2984 259420 2990
rect 259368 2926 259420 2932
rect 258276 480 258304 2926
rect 259472 480 259500 3334
rect 260668 480 260696 4966
rect 261772 480 261800 9998
rect 263336 6914 263364 49030
rect 263428 26926 263456 87774
rect 264348 85542 264376 87774
rect 265268 85542 265296 87774
rect 263508 85536 263560 85542
rect 263508 85478 263560 85484
rect 264336 85536 264388 85542
rect 264336 85478 264388 85484
rect 264888 85536 264940 85542
rect 264888 85478 264940 85484
rect 265256 85536 265308 85542
rect 265256 85478 265308 85484
rect 263416 26920 263468 26926
rect 263416 26862 263468 26868
rect 263520 24138 263548 85478
rect 264900 29646 264928 85478
rect 264888 29640 264940 29646
rect 264888 29582 264940 29588
rect 263508 24132 263560 24138
rect 263508 24074 263560 24080
rect 266084 9988 266136 9994
rect 266084 9930 266136 9936
rect 262968 6886 263364 6914
rect 262968 480 262996 6886
rect 264152 4820 264204 4826
rect 264152 4762 264204 4768
rect 264164 480 264192 4762
rect 266096 3398 266124 9930
rect 266188 4826 266216 87774
rect 267108 85542 267136 87774
rect 268028 85542 268056 87774
rect 266268 85536 266320 85542
rect 266268 85478 266320 85484
rect 267096 85536 267148 85542
rect 267096 85478 267148 85484
rect 267648 85536 267700 85542
rect 267648 85478 267700 85484
rect 268016 85536 268068 85542
rect 268016 85478 268068 85484
rect 266280 5030 266308 85478
rect 267004 85332 267056 85338
rect 267004 85274 267056 85280
rect 267016 21418 267044 85274
rect 267556 51808 267608 51814
rect 267556 51750 267608 51756
rect 267004 21412 267056 21418
rect 267004 21354 267056 21360
rect 266268 5024 266320 5030
rect 266268 4966 266320 4972
rect 266176 4820 266228 4826
rect 266176 4762 266228 4768
rect 267568 3398 267596 51750
rect 267660 4214 267688 85478
rect 268844 9920 268896 9926
rect 268844 9862 268896 9868
rect 267740 5296 267792 5302
rect 267740 5238 267792 5244
rect 267648 4208 267700 4214
rect 267648 4150 267700 4156
rect 265348 3392 265400 3398
rect 265348 3334 265400 3340
rect 266084 3392 266136 3398
rect 266084 3334 266136 3340
rect 266544 3392 266596 3398
rect 266544 3334 266596 3340
rect 267556 3392 267608 3398
rect 267556 3334 267608 3340
rect 265360 480 265388 3334
rect 266556 480 266584 3334
rect 267752 480 267780 5238
rect 268856 480 268884 9862
rect 268948 4486 268976 87774
rect 269868 85542 269896 87774
rect 270788 85542 270816 87774
rect 269028 85536 269080 85542
rect 269028 85478 269080 85484
rect 269856 85536 269908 85542
rect 269856 85478 269908 85484
rect 270408 85536 270460 85542
rect 270408 85478 270460 85484
rect 270776 85536 270828 85542
rect 270776 85478 270828 85484
rect 268936 4480 268988 4486
rect 268936 4422 268988 4428
rect 269040 4282 269068 85478
rect 270040 11076 270092 11082
rect 270040 11018 270092 11024
rect 269028 4276 269080 4282
rect 269028 4218 269080 4224
rect 270052 480 270080 11018
rect 270420 4554 270448 85478
rect 271616 84194 271644 87774
rect 272536 85542 272564 87774
rect 273456 85542 273484 87774
rect 271788 85536 271840 85542
rect 271788 85478 271840 85484
rect 272524 85536 272576 85542
rect 272524 85478 272576 85484
rect 273168 85536 273220 85542
rect 273168 85478 273220 85484
rect 273444 85536 273496 85542
rect 273444 85478 273496 85484
rect 271616 84166 271736 84194
rect 271236 5228 271288 5234
rect 271236 5170 271288 5176
rect 270408 4548 270460 4554
rect 270408 4490 270460 4496
rect 271248 480 271276 5170
rect 271708 4758 271736 84166
rect 271800 5234 271828 85478
rect 273076 9716 273128 9722
rect 273076 9658 273128 9664
rect 271788 5228 271840 5234
rect 271788 5170 271840 5176
rect 271696 4752 271748 4758
rect 271696 4694 271748 4700
rect 273088 3398 273116 9658
rect 273180 4622 273208 85478
rect 274376 84194 274404 87774
rect 275296 85542 275324 87774
rect 276216 85542 276244 87774
rect 277136 86954 277164 87774
rect 277136 86926 277348 86954
rect 274548 85536 274600 85542
rect 274548 85478 274600 85484
rect 275284 85536 275336 85542
rect 275284 85478 275336 85484
rect 275928 85536 275980 85542
rect 275928 85478 275980 85484
rect 276204 85536 276256 85542
rect 276204 85478 276256 85484
rect 277216 85536 277268 85542
rect 277216 85478 277268 85484
rect 274376 84166 274496 84194
rect 274364 73840 274416 73846
rect 274364 73782 274416 73788
rect 273258 9072 273314 9081
rect 273258 9007 273314 9016
rect 273272 8974 273300 9007
rect 273260 8968 273312 8974
rect 273352 8968 273404 8974
rect 273260 8910 273312 8916
rect 273350 8936 273352 8945
rect 273404 8936 273406 8945
rect 273350 8871 273406 8880
rect 273168 4616 273220 4622
rect 273168 4558 273220 4564
rect 274376 4146 274404 73782
rect 274468 5370 274496 84166
rect 274456 5364 274508 5370
rect 274456 5306 274508 5312
rect 274560 5302 274588 85478
rect 275940 5574 275968 85478
rect 277228 12434 277256 85478
rect 277136 12406 277256 12434
rect 275928 5568 275980 5574
rect 275928 5510 275980 5516
rect 277136 5370 277164 12406
rect 277320 10554 277348 86926
rect 278056 85542 278084 87774
rect 278976 85542 279004 87774
rect 278044 85536 278096 85542
rect 278044 85478 278096 85484
rect 278688 85536 278740 85542
rect 278688 85478 278740 85484
rect 278964 85536 279016 85542
rect 278964 85478 279016 85484
rect 278044 58676 278096 58682
rect 278044 58618 278096 58624
rect 277228 10526 277348 10554
rect 277124 5364 277176 5370
rect 277124 5306 277176 5312
rect 274548 5296 274600 5302
rect 274548 5238 274600 5244
rect 277228 5166 277256 10526
rect 277306 10432 277362 10441
rect 277306 10367 277362 10376
rect 274824 5160 274876 5166
rect 274824 5102 274876 5108
rect 277216 5160 277268 5166
rect 277216 5102 277268 5108
rect 273628 4140 273680 4146
rect 273628 4082 273680 4088
rect 274364 4140 274416 4146
rect 274364 4082 274416 4088
rect 272432 3392 272484 3398
rect 272432 3334 272484 3340
rect 273076 3392 273128 3398
rect 273076 3334 273128 3340
rect 272444 480 272472 3334
rect 273640 480 273668 4082
rect 274836 480 274864 5102
rect 277216 4140 277268 4146
rect 277216 4082 277268 4088
rect 276020 3936 276072 3942
rect 276020 3878 276072 3884
rect 276032 480 276060 3878
rect 277228 1986 277256 4082
rect 277320 3942 277348 10367
rect 278056 4146 278084 58618
rect 278700 5370 278728 85478
rect 279804 85338 279832 87774
rect 280724 85542 280752 87774
rect 280068 85536 280120 85542
rect 280068 85478 280120 85484
rect 280160 85536 280212 85542
rect 280160 85478 280212 85484
rect 280712 85536 280764 85542
rect 280712 85478 280764 85484
rect 280804 85536 280856 85542
rect 280804 85478 280856 85484
rect 279792 85332 279844 85338
rect 279792 85274 279844 85280
rect 279514 10160 279570 10169
rect 279514 10095 279570 10104
rect 278688 5364 278740 5370
rect 278688 5306 278740 5312
rect 278320 5092 278372 5098
rect 278320 5034 278372 5040
rect 278044 4140 278096 4146
rect 278044 4082 278096 4088
rect 277308 3936 277360 3942
rect 277308 3878 277360 3884
rect 277136 1958 277256 1986
rect 277136 480 277164 1958
rect 278332 480 278360 5034
rect 279528 480 279556 10095
rect 280080 4078 280108 85478
rect 280172 77994 280200 85478
rect 280160 77988 280212 77994
rect 280160 77930 280212 77936
rect 280816 24274 280844 85478
rect 281644 85338 281672 87774
rect 282564 85542 282592 87774
rect 283392 87774 283500 87802
rect 284312 87774 284420 87802
rect 285232 87774 285340 87802
rect 286232 87802 286260 88049
rect 287060 87802 287088 88049
rect 287980 87802 288008 88049
rect 288900 87802 288928 88049
rect 286232 87774 286272 87802
rect 287060 87774 287100 87802
rect 282552 85536 282604 85542
rect 282552 85478 282604 85484
rect 280896 85332 280948 85338
rect 280896 85274 280948 85280
rect 281632 85332 281684 85338
rect 281632 85274 281684 85280
rect 280908 75206 280936 85274
rect 283392 84194 283420 87774
rect 282932 84166 283420 84194
rect 281448 76560 281500 76566
rect 281448 76502 281500 76508
rect 280896 75200 280948 75206
rect 280896 75142 280948 75148
rect 280804 24268 280856 24274
rect 280804 24210 280856 24216
rect 280068 4072 280120 4078
rect 280068 4014 280120 4020
rect 281460 2922 281488 76502
rect 281540 32564 281592 32570
rect 281540 32506 281592 32512
rect 281552 16574 281580 32506
rect 281552 16546 281948 16574
rect 280712 2916 280764 2922
rect 280712 2858 280764 2864
rect 281448 2916 281500 2922
rect 281448 2858 281500 2864
rect 280724 480 280752 2858
rect 281920 480 281948 16546
rect 282644 11076 282696 11082
rect 282644 11018 282696 11024
rect 282656 10985 282684 11018
rect 282642 10976 282698 10985
rect 282642 10911 282698 10920
rect 282828 10464 282880 10470
rect 282826 10432 282828 10441
rect 282880 10432 282882 10441
rect 282826 10367 282882 10376
rect 282932 9081 282960 84166
rect 284312 35222 284340 87774
rect 285232 84194 285260 87774
rect 286244 84998 286272 87774
rect 286416 85332 286468 85338
rect 286416 85274 286468 85280
rect 286232 84992 286284 84998
rect 286232 84934 286284 84940
rect 284404 84166 285260 84194
rect 286324 84244 286376 84250
rect 286324 84186 286376 84192
rect 284404 78062 284432 84166
rect 284392 78056 284444 78062
rect 284392 77998 284444 78004
rect 285588 53168 285640 53174
rect 285588 53110 285640 53116
rect 284484 35488 284536 35494
rect 284484 35430 284536 35436
rect 284300 35216 284352 35222
rect 284300 35158 284352 35164
rect 284496 16574 284524 35430
rect 284496 16546 285444 16574
rect 282918 9072 282974 9081
rect 282918 9007 282974 9016
rect 284208 7404 284260 7410
rect 284208 7346 284260 7352
rect 282828 5636 282880 5642
rect 282828 5578 282880 5584
rect 282840 5302 282868 5578
rect 282828 5296 282880 5302
rect 282828 5238 282880 5244
rect 284220 4146 284248 7346
rect 283104 4140 283156 4146
rect 283104 4082 283156 4088
rect 284208 4140 284260 4146
rect 284208 4082 284260 4088
rect 284300 4140 284352 4146
rect 284300 4082 284352 4088
rect 283116 480 283144 4082
rect 284312 480 284340 4082
rect 285416 480 285444 16546
rect 285600 4146 285628 53110
rect 286336 29714 286364 84186
rect 286428 35222 286456 85274
rect 287072 84250 287100 87774
rect 287624 87774 288008 87802
rect 288820 87774 288928 87802
rect 289820 87802 289848 88049
rect 290740 87802 290768 88049
rect 291660 87802 291688 88049
rect 289820 87774 289860 87802
rect 287060 84244 287112 84250
rect 287624 84194 287652 87774
rect 287704 84992 287756 84998
rect 287704 84934 287756 84940
rect 287060 84186 287112 84192
rect 287164 84166 287652 84194
rect 287164 73914 287192 84166
rect 287152 73908 287204 73914
rect 287152 73850 287204 73856
rect 286416 35216 286468 35222
rect 286416 35158 286468 35164
rect 286324 29708 286376 29714
rect 286324 29650 286376 29656
rect 287716 14618 287744 84934
rect 288820 84194 288848 87774
rect 289832 85542 289860 87774
rect 290660 87774 290768 87802
rect 291580 87774 291688 87802
rect 292580 87802 292608 88049
rect 293500 87802 293528 88049
rect 294328 87802 294356 88049
rect 292580 87774 292620 87802
rect 289084 85536 289136 85542
rect 289084 85478 289136 85484
rect 289820 85536 289872 85542
rect 289820 85478 289872 85484
rect 288452 84166 288848 84194
rect 288452 83570 288480 84166
rect 288440 83564 288492 83570
rect 288440 83506 288492 83512
rect 289096 75274 289124 85478
rect 290660 84194 290688 87774
rect 291580 84194 291608 87774
rect 289924 84166 290688 84194
rect 291212 84166 291608 84194
rect 289084 75268 289136 75274
rect 289084 75210 289136 75216
rect 288440 38208 288492 38214
rect 288440 38150 288492 38156
rect 288348 35284 288400 35290
rect 288348 35226 288400 35232
rect 287704 14612 287756 14618
rect 287704 14554 287756 14560
rect 286600 6724 286652 6730
rect 286600 6666 286652 6672
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 286612 480 286640 6666
rect 288360 4146 288388 35226
rect 288452 16574 288480 38150
rect 289924 18766 289952 84166
rect 291212 26994 291240 84166
rect 292488 83564 292540 83570
rect 292488 83506 292540 83512
rect 291200 26988 291252 26994
rect 291200 26930 291252 26936
rect 289912 18760 289964 18766
rect 289912 18702 289964 18708
rect 288452 16546 289032 16574
rect 287796 4140 287848 4146
rect 287796 4082 287848 4088
rect 288348 4140 288400 4146
rect 288348 4082 288400 4088
rect 287808 480 287836 4082
rect 289004 480 289032 16546
rect 292304 11144 292356 11150
rect 292302 11112 292304 11121
rect 292356 11112 292358 11121
rect 292302 11047 292358 11056
rect 292396 10532 292448 10538
rect 292396 10474 292448 10480
rect 292408 10169 292436 10474
rect 292394 10160 292450 10169
rect 292394 10095 292450 10104
rect 292396 9512 292448 9518
rect 292396 9454 292448 9460
rect 292408 9353 292436 9454
rect 292394 9344 292450 9353
rect 292394 9279 292450 9288
rect 290188 6792 290240 6798
rect 290188 6734 290240 6740
rect 290200 480 290228 6734
rect 292500 4146 292528 83506
rect 292592 11257 292620 87774
rect 293420 87774 293528 87802
rect 294248 87774 294356 87802
rect 295248 87802 295276 88049
rect 296168 87802 296196 88049
rect 295248 87774 295288 87802
rect 293420 84194 293448 87774
rect 294248 86954 294276 87774
rect 292684 84166 293448 84194
rect 293972 86926 294276 86954
rect 292578 11248 292634 11257
rect 292578 11183 292634 11192
rect 292580 11076 292632 11082
rect 292580 11018 292632 11024
rect 292592 10849 292620 11018
rect 292578 10840 292634 10849
rect 292578 10775 292634 10784
rect 292684 9382 292712 84166
rect 292764 17332 292816 17338
rect 292764 17274 292816 17280
rect 292672 9376 292724 9382
rect 292672 9318 292724 9324
rect 291384 4140 291436 4146
rect 291384 4082 291436 4088
rect 292488 4140 292540 4146
rect 292488 4082 292540 4088
rect 291396 480 291424 4082
rect 292776 2774 292804 17274
rect 292854 11248 292910 11257
rect 292854 11183 292910 11192
rect 292868 9110 292896 11183
rect 292948 11144 293000 11150
rect 292946 11112 292948 11121
rect 293000 11112 293002 11121
rect 292946 11047 293002 11056
rect 293972 9518 294000 86926
rect 295260 86154 295288 87774
rect 296088 87774 296196 87802
rect 296720 87848 296772 87854
rect 297088 87802 297116 88049
rect 298008 87854 298036 88049
rect 296720 87790 296772 87796
rect 294052 86148 294104 86154
rect 294052 86090 294104 86096
rect 295248 86148 295300 86154
rect 295248 86090 295300 86096
rect 293960 9512 294012 9518
rect 293960 9454 294012 9460
rect 294064 9450 294092 86090
rect 296088 84194 296116 87774
rect 295352 84166 296116 84194
rect 295248 26988 295300 26994
rect 295248 26930 295300 26936
rect 294052 9444 294104 9450
rect 294052 9386 294104 9392
rect 292948 9376 293000 9382
rect 292946 9344 292948 9353
rect 293000 9344 293002 9353
rect 292946 9279 293002 9288
rect 292856 9104 292908 9110
rect 292856 9046 292908 9052
rect 293684 6860 293736 6866
rect 293684 6802 293736 6808
rect 292592 2746 292804 2774
rect 292592 480 292620 2746
rect 293696 480 293724 6802
rect 295260 2774 295288 26930
rect 295352 9382 295380 84166
rect 295432 39432 295484 39438
rect 295432 39374 295484 39380
rect 295444 16574 295472 39374
rect 295444 16546 296116 16574
rect 295340 9376 295392 9382
rect 295340 9318 295392 9324
rect 294892 2746 295288 2774
rect 294892 480 294920 2746
rect 296088 480 296116 16546
rect 296732 9586 296760 87790
rect 297008 87774 297116 87802
rect 297996 87848 298048 87854
rect 298928 87802 298956 88049
rect 297996 87790 298048 87796
rect 298848 87774 298956 87802
rect 299480 87848 299532 87854
rect 299848 87802 299876 88049
rect 300768 87854 300796 88049
rect 299480 87790 299532 87796
rect 297008 84194 297036 87774
rect 298848 84194 298876 87774
rect 296824 84166 297036 84194
rect 298112 84166 298876 84194
rect 296824 16574 296852 84166
rect 296824 16546 297036 16574
rect 296720 9580 296772 9586
rect 296720 9522 296772 9528
rect 297008 9178 297036 16546
rect 298112 9654 298140 84166
rect 299388 55956 299440 55962
rect 299388 55898 299440 55904
rect 298100 9648 298152 9654
rect 298100 9590 298152 9596
rect 296996 9172 297048 9178
rect 296996 9114 297048 9120
rect 297272 6112 297324 6118
rect 297272 6054 297324 6060
rect 297284 480 297312 6054
rect 299400 4146 299428 55898
rect 299492 8838 299520 87790
rect 299768 87774 299876 87802
rect 300756 87848 300808 87854
rect 301596 87802 301624 88049
rect 302516 87802 302544 88049
rect 303436 87802 303464 88049
rect 304356 87802 304384 88049
rect 305276 87802 305304 88049
rect 306196 87802 306224 88049
rect 307116 87802 307144 88049
rect 308036 87802 308064 88049
rect 308864 87802 308892 88049
rect 300756 87790 300808 87796
rect 301516 87774 301624 87802
rect 302252 87774 302544 87802
rect 303356 87774 303464 87802
rect 304276 87774 304384 87802
rect 305012 87774 305304 87802
rect 306116 87774 306224 87802
rect 307036 87774 307144 87802
rect 307956 87774 308064 87802
rect 308324 87774 308892 87802
rect 309784 87802 309812 88049
rect 310704 87802 310732 88049
rect 311624 87802 311652 88049
rect 312544 87802 312572 88049
rect 309784 87774 309824 87802
rect 310704 87774 310744 87802
rect 311624 87774 311664 87802
rect 299768 84194 299796 87774
rect 301516 84194 301544 87774
rect 299584 84166 299796 84194
rect 300872 84166 301544 84194
rect 299584 8906 299612 84166
rect 299664 42152 299716 42158
rect 299664 42094 299716 42100
rect 299572 8900 299624 8906
rect 299572 8842 299624 8848
rect 299480 8832 299532 8838
rect 299480 8774 299532 8780
rect 298468 4140 298520 4146
rect 298468 4082 298520 4088
rect 299388 4140 299440 4146
rect 299388 4082 299440 4088
rect 298480 480 298508 4082
rect 299676 480 299704 42094
rect 300872 8634 300900 84166
rect 302148 22772 302200 22778
rect 302148 22714 302200 22720
rect 300860 8628 300912 8634
rect 300860 8570 300912 8576
rect 300768 5908 300820 5914
rect 300768 5850 300820 5856
rect 300780 480 300808 5850
rect 302160 2774 302188 22714
rect 302252 8566 302280 87774
rect 303356 84194 303384 87774
rect 304276 84194 304304 87774
rect 302344 84166 303384 84194
rect 303632 84166 304304 84194
rect 302344 12434 302372 84166
rect 302424 44940 302476 44946
rect 302424 44882 302476 44888
rect 302436 16574 302464 44882
rect 302436 16546 303200 16574
rect 302344 12406 302464 12434
rect 302330 10840 302386 10849
rect 302330 10775 302332 10784
rect 302384 10775 302386 10784
rect 302332 10746 302384 10752
rect 302332 10532 302384 10538
rect 302332 10474 302384 10480
rect 302344 10169 302372 10474
rect 302330 10160 302386 10169
rect 302330 10095 302386 10104
rect 302240 8560 302292 8566
rect 302240 8502 302292 8508
rect 302436 8498 302464 12406
rect 302514 11112 302570 11121
rect 302514 11047 302516 11056
rect 302568 11047 302570 11056
rect 302516 11018 302568 11024
rect 302424 8492 302476 8498
rect 302424 8434 302476 8440
rect 301976 2746 302188 2774
rect 301976 480 302004 2746
rect 303172 480 303200 16546
rect 303632 8430 303660 84166
rect 303620 8424 303672 8430
rect 303620 8366 303672 8372
rect 305012 8362 305040 87774
rect 306116 84194 306144 87774
rect 307036 84194 307064 87774
rect 307956 86954 307984 87774
rect 305104 84166 306144 84194
rect 306392 84166 307064 84194
rect 307772 86926 307984 86954
rect 305104 8974 305132 84166
rect 306392 29782 306420 84166
rect 307772 75342 307800 86926
rect 308324 84194 308352 87774
rect 309796 85542 309824 87774
rect 310716 85542 310744 87774
rect 308404 85536 308456 85542
rect 308404 85478 308456 85484
rect 309784 85536 309836 85542
rect 309784 85478 309836 85484
rect 309876 85536 309928 85542
rect 309876 85478 309928 85484
rect 310704 85536 310756 85542
rect 310704 85478 310756 85484
rect 307864 84166 308352 84194
rect 307864 78130 307892 84166
rect 307852 78124 307904 78130
rect 307852 78066 307904 78072
rect 307760 75336 307812 75342
rect 307760 75278 307812 75284
rect 306472 47660 306524 47666
rect 306472 47602 306524 47608
rect 306380 29776 306432 29782
rect 306380 29718 306432 29724
rect 306484 16574 306512 47602
rect 308416 22982 308444 85478
rect 309784 82272 309836 82278
rect 309784 82214 309836 82220
rect 308496 57316 308548 57322
rect 308496 57258 308548 57264
rect 308404 22976 308456 22982
rect 308404 22918 308456 22924
rect 306484 16546 306788 16574
rect 305092 8968 305144 8974
rect 305092 8910 305144 8916
rect 305000 8356 305052 8362
rect 305000 8298 305052 8304
rect 304356 5840 304408 5846
rect 304356 5782 304408 5788
rect 304368 480 304396 5782
rect 305552 4140 305604 4146
rect 305552 4082 305604 4088
rect 305564 480 305592 4082
rect 306760 480 306788 16546
rect 307944 5772 307996 5778
rect 307944 5714 307996 5720
rect 307956 480 307984 5714
rect 308508 4146 308536 57258
rect 309140 50448 309192 50454
rect 309140 50390 309192 50396
rect 309152 16574 309180 50390
rect 309152 16546 309732 16574
rect 308496 4140 308548 4146
rect 308496 4082 308548 4088
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 309060 480 309088 4082
rect 309704 2774 309732 16546
rect 309796 4146 309824 82214
rect 309888 31142 309916 85478
rect 311636 85338 311664 87774
rect 312464 87774 312572 87802
rect 313464 87802 313492 88049
rect 314384 87802 314412 88049
rect 315304 87802 315332 88049
rect 313464 87774 313504 87802
rect 310428 85332 310480 85338
rect 310428 85274 310480 85280
rect 311624 85332 311676 85338
rect 311624 85274 311676 85280
rect 310440 80850 310468 85274
rect 312464 84194 312492 87774
rect 313476 85542 313504 87774
rect 314304 87774 314412 87802
rect 315224 87774 315332 87802
rect 316040 87848 316092 87854
rect 316040 87790 316092 87796
rect 316132 87802 316160 88049
rect 317052 87854 317080 88049
rect 317040 87848 317092 87854
rect 312544 85536 312596 85542
rect 312544 85478 312596 85484
rect 313464 85536 313516 85542
rect 313464 85478 313516 85484
rect 311912 84166 312492 84194
rect 310428 80844 310480 80850
rect 310428 80786 310480 80792
rect 309876 31136 309928 31142
rect 309876 31078 309928 31084
rect 311912 25702 311940 84166
rect 312556 28422 312584 85478
rect 314304 84194 314332 87774
rect 315224 84194 315252 87774
rect 313476 84166 314332 84194
rect 314672 84166 315252 84194
rect 313372 53236 313424 53242
rect 313372 53178 313424 53184
rect 312544 28416 312596 28422
rect 312544 28358 312596 28364
rect 311900 25696 311952 25702
rect 311900 25638 311952 25644
rect 313188 25696 313240 25702
rect 313188 25638 313240 25644
rect 311808 10736 311860 10742
rect 311636 10684 311808 10690
rect 311636 10678 311860 10684
rect 311636 10662 311848 10678
rect 311532 10464 311584 10470
rect 311438 10432 311494 10441
rect 311532 10406 311584 10412
rect 311438 10367 311494 10376
rect 311452 10266 311480 10367
rect 311440 10260 311492 10266
rect 311440 10202 311492 10208
rect 311544 10010 311572 10406
rect 311636 10198 311664 10662
rect 311808 10260 311860 10266
rect 311808 10202 311860 10208
rect 311624 10192 311676 10198
rect 311716 10192 311768 10198
rect 311624 10134 311676 10140
rect 311714 10160 311716 10169
rect 311768 10160 311770 10169
rect 311714 10095 311770 10104
rect 311820 10010 311848 10202
rect 311544 9982 311848 10010
rect 311440 5636 311492 5642
rect 311440 5578 311492 5584
rect 309784 4140 309836 4146
rect 309784 4082 309836 4088
rect 309704 2746 310284 2774
rect 310256 480 310284 2746
rect 311452 480 311480 5578
rect 313200 3398 313228 25638
rect 313384 6914 313412 53178
rect 313476 10441 313504 84166
rect 313462 10432 313518 10441
rect 313462 10367 313518 10376
rect 314672 9654 314700 84166
rect 316052 9994 316080 87790
rect 316132 87774 316172 87802
rect 317972 87802 318000 88049
rect 318892 87802 318920 88049
rect 319812 87802 319840 88049
rect 320732 87802 320760 88049
rect 317040 87790 317092 87796
rect 316144 10130 316172 87774
rect 317892 87774 318000 87802
rect 318812 87774 318920 87802
rect 319732 87774 319840 87802
rect 320652 87774 320760 87802
rect 321560 87848 321612 87854
rect 321560 87790 321612 87796
rect 321652 87802 321680 88049
rect 322572 87854 322600 88049
rect 322560 87848 322612 87854
rect 317892 84194 317920 87774
rect 317432 84166 317920 84194
rect 316224 56160 316276 56166
rect 316224 56102 316276 56108
rect 316236 16574 316264 56102
rect 316236 16546 317368 16574
rect 316132 10124 316184 10130
rect 316132 10066 316184 10072
rect 316040 9988 316092 9994
rect 316040 9930 316092 9936
rect 314660 9648 314712 9654
rect 314660 9590 314712 9596
rect 313384 6886 313872 6914
rect 312636 3392 312688 3398
rect 312636 3334 312688 3340
rect 313188 3392 313240 3398
rect 313188 3334 313240 3340
rect 312648 480 312676 3334
rect 313844 480 313872 6886
rect 315028 5704 315080 5710
rect 315028 5646 315080 5652
rect 315040 480 315068 5646
rect 316040 5568 316092 5574
rect 316040 5510 316092 5516
rect 316052 5001 316080 5510
rect 316038 4992 316094 5001
rect 316038 4927 316094 4936
rect 316224 3392 316276 3398
rect 316224 3334 316276 3340
rect 316236 480 316264 3334
rect 317340 480 317368 16546
rect 317432 10062 317460 84166
rect 318064 60104 318116 60110
rect 318064 60046 318116 60052
rect 317420 10056 317472 10062
rect 317420 9998 317472 10004
rect 318076 3398 318104 60046
rect 318812 9926 318840 87774
rect 319732 84194 319760 87774
rect 320652 84194 320680 87774
rect 318904 84166 319760 84194
rect 320192 84166 320680 84194
rect 318800 9920 318852 9926
rect 318800 9862 318852 9868
rect 318904 9722 318932 84166
rect 320192 10266 320220 84166
rect 320272 57384 320324 57390
rect 320272 57326 320324 57332
rect 320284 16574 320312 57326
rect 320824 28416 320876 28422
rect 320824 28358 320876 28364
rect 320284 16546 320772 16574
rect 320180 10260 320232 10266
rect 320180 10202 320232 10208
rect 318892 9716 318944 9722
rect 318892 9658 318944 9664
rect 318524 5568 318576 5574
rect 318524 5510 318576 5516
rect 318064 3392 318116 3398
rect 318064 3334 318116 3340
rect 318536 480 318564 5510
rect 319720 3732 319772 3738
rect 319720 3674 319772 3680
rect 319732 480 319760 3674
rect 320744 3482 320772 16546
rect 320836 3738 320864 28358
rect 321572 9042 321600 87790
rect 321652 87774 321692 87802
rect 323400 87802 323428 88049
rect 322560 87790 322612 87796
rect 321664 10198 321692 87774
rect 323320 87774 323428 87802
rect 324320 87802 324348 88049
rect 325240 87802 325268 88049
rect 326160 87802 326188 88049
rect 324320 87774 324360 87802
rect 323320 84194 323348 87774
rect 322952 84166 323348 84194
rect 321652 10192 321704 10198
rect 321652 10134 321704 10140
rect 321560 9036 321612 9042
rect 321560 8978 321612 8984
rect 322952 6730 322980 84166
rect 324228 62892 324280 62898
rect 324228 62834 324280 62840
rect 322940 6724 322992 6730
rect 322940 6666 322992 6672
rect 323032 6724 323084 6730
rect 323032 6666 323084 6672
rect 323044 6610 323072 6666
rect 322860 6582 323072 6610
rect 320824 3732 320876 3738
rect 320824 3674 320876 3680
rect 320744 3454 320956 3482
rect 320928 480 320956 3454
rect 322860 3194 322888 6582
rect 324240 3398 324268 62834
rect 324332 6798 324360 87774
rect 325160 87774 325268 87802
rect 326080 87774 326188 87802
rect 327080 87802 327108 88049
rect 328000 87802 328028 88049
rect 328920 87802 328948 88049
rect 327080 87774 327120 87802
rect 325160 84194 325188 87774
rect 326080 84194 326108 87774
rect 324424 84166 325188 84194
rect 325712 84166 326108 84194
rect 324424 6866 324452 84166
rect 324504 60172 324556 60178
rect 324504 60114 324556 60120
rect 324412 6860 324464 6866
rect 324412 6802 324464 6808
rect 324320 6792 324372 6798
rect 324320 6734 324372 6740
rect 324516 3482 324544 60114
rect 325608 6792 325660 6798
rect 325608 6734 325660 6740
rect 324424 3454 324544 3482
rect 323308 3392 323360 3398
rect 323308 3334 323360 3340
rect 324228 3392 324280 3398
rect 324228 3334 324280 3340
rect 322112 3188 322164 3194
rect 322112 3130 322164 3136
rect 322848 3188 322900 3194
rect 322848 3130 322900 3136
rect 322124 480 322152 3130
rect 323320 480 323348 3334
rect 324424 480 324452 3454
rect 325620 480 325648 6734
rect 325712 6118 325740 84166
rect 326988 29708 327040 29714
rect 326988 29650 327040 29656
rect 327000 6914 327028 29650
rect 326816 6886 327028 6914
rect 325700 6112 325752 6118
rect 325700 6054 325752 6060
rect 326816 480 326844 6886
rect 327092 5914 327120 87774
rect 327920 87774 328028 87802
rect 328840 87774 328948 87802
rect 329840 87802 329868 88049
rect 330668 87802 330696 88049
rect 331588 87802 331616 88049
rect 329840 87774 329880 87802
rect 327920 84194 327948 87774
rect 328840 84194 328868 87774
rect 327184 84166 327948 84194
rect 328472 84166 328868 84194
rect 327080 5908 327132 5914
rect 327080 5850 327132 5856
rect 327184 5846 327212 84166
rect 327264 62960 327316 62966
rect 327264 62902 327316 62908
rect 327276 16574 327304 62902
rect 327276 16546 328040 16574
rect 327172 5840 327224 5846
rect 327172 5782 327224 5788
rect 328012 480 328040 16546
rect 328472 5778 328500 84166
rect 328460 5772 328512 5778
rect 328460 5714 328512 5720
rect 329852 5710 329880 87774
rect 330588 87774 330696 87802
rect 331508 87774 331616 87802
rect 332508 87802 332536 88049
rect 333428 87802 333456 88049
rect 332508 87774 332548 87802
rect 330588 84194 330616 87774
rect 331508 87258 331536 87774
rect 329944 84166 330616 84194
rect 331232 87230 331536 87258
rect 329840 5704 329892 5710
rect 329840 5646 329892 5652
rect 329196 5636 329248 5642
rect 329196 5578 329248 5584
rect 329208 480 329236 5578
rect 329944 5574 329972 84166
rect 331128 31136 331180 31142
rect 331128 31078 331180 31084
rect 329932 5568 329984 5574
rect 329932 5510 329984 5516
rect 331140 3398 331168 31078
rect 331232 5846 331260 87230
rect 332520 86154 332548 87774
rect 333348 87774 333456 87802
rect 333980 87848 334032 87854
rect 334348 87802 334376 88049
rect 335268 87854 335296 88049
rect 333980 87790 334032 87796
rect 331312 86148 331364 86154
rect 331312 86090 331364 86096
rect 332508 86148 332560 86154
rect 332508 86090 332560 86096
rect 331324 6730 331352 86090
rect 333348 84194 333376 87774
rect 332612 84166 333376 84194
rect 331404 65612 331456 65618
rect 331404 65554 331456 65560
rect 331416 16574 331444 65554
rect 331416 16546 331628 16574
rect 331312 6724 331364 6730
rect 331312 6666 331364 6672
rect 331220 5840 331272 5846
rect 331220 5782 331272 5788
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 331128 3392 331180 3398
rect 331128 3334 331180 3340
rect 330404 480 330432 3334
rect 331600 480 331628 16546
rect 332612 6798 332640 84166
rect 332600 6792 332652 6798
rect 332600 6734 332652 6740
rect 333992 5574 334020 87790
rect 334268 87774 334376 87802
rect 335256 87848 335308 87854
rect 336188 87802 336216 88049
rect 335256 87790 335308 87796
rect 336108 87774 336216 87802
rect 337108 87802 337136 88049
rect 337936 87802 337964 88049
rect 338856 87802 338884 88049
rect 339776 87802 339804 88049
rect 340696 87802 340724 88049
rect 341616 87802 341644 88049
rect 342536 87802 342564 88049
rect 343456 87802 343484 88049
rect 344376 87802 344404 88049
rect 345204 87802 345232 88049
rect 346124 87802 346152 88049
rect 347044 87802 347072 88049
rect 347964 87802 347992 88049
rect 348884 87802 348912 88049
rect 349804 87802 349832 88049
rect 350724 87802 350752 88049
rect 351644 87802 351672 88049
rect 352472 87802 352500 88049
rect 353392 87802 353420 88049
rect 354312 87938 354340 88049
rect 354312 87910 354628 87938
rect 337108 87774 337148 87802
rect 337936 87774 337976 87802
rect 338856 87774 338896 87802
rect 339776 87774 339816 87802
rect 340696 87774 340736 87802
rect 341616 87774 341656 87802
rect 342536 87774 342576 87802
rect 343456 87774 343588 87802
rect 344376 87774 344416 87802
rect 345204 87774 345244 87802
rect 346124 87774 346164 87802
rect 347044 87774 347084 87802
rect 347964 87774 348004 87802
rect 348884 87774 348924 87802
rect 349804 87774 349844 87802
rect 350724 87774 350764 87802
rect 351644 87774 351684 87802
rect 352472 87774 352512 87802
rect 353392 87774 353432 87802
rect 334268 84194 334296 87774
rect 336108 84194 336136 87774
rect 337120 85542 337148 87774
rect 337108 85536 337160 85542
rect 337108 85478 337160 85484
rect 334084 84166 334296 84194
rect 335372 84166 336136 84194
rect 334084 5642 334112 84166
rect 334164 68400 334216 68406
rect 334164 68342 334216 68348
rect 334176 16574 334204 68342
rect 334176 16546 335124 16574
rect 334072 5636 334124 5642
rect 334072 5578 334124 5584
rect 334164 5636 334216 5642
rect 334164 5578 334216 5584
rect 332692 5568 332744 5574
rect 332692 5510 332744 5516
rect 333980 5568 334032 5574
rect 333980 5510 334032 5516
rect 332704 480 332732 5510
rect 334176 5001 334204 5578
rect 334162 4992 334218 5001
rect 334162 4927 334218 4936
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 333900 480 333928 3946
rect 335096 480 335124 16546
rect 335372 3398 335400 84166
rect 336004 39432 336056 39438
rect 336004 39374 336056 39380
rect 336016 4010 336044 39374
rect 337948 5846 337976 87774
rect 338868 85542 338896 87774
rect 339788 85542 339816 87774
rect 338028 85536 338080 85542
rect 338028 85478 338080 85484
rect 338856 85536 338908 85542
rect 338856 85478 338908 85484
rect 339408 85536 339460 85542
rect 339408 85478 339460 85484
rect 339776 85536 339828 85542
rect 339776 85478 339828 85484
rect 337936 5840 337988 5846
rect 337936 5782 337988 5788
rect 338040 5642 338068 85478
rect 338120 71120 338172 71126
rect 338120 71062 338172 71068
rect 338132 16574 338160 71062
rect 338764 42220 338816 42226
rect 338764 42162 338816 42168
rect 338132 16546 338712 16574
rect 338028 5636 338080 5642
rect 338028 5578 338080 5584
rect 336004 4004 336056 4010
rect 336004 3946 336056 3952
rect 335360 3392 335412 3398
rect 335360 3334 335412 3340
rect 336280 3392 336332 3398
rect 336280 3334 336332 3340
rect 337476 3392 337528 3398
rect 337476 3334 337528 3340
rect 336292 480 336320 3334
rect 337488 480 337516 3334
rect 338684 480 338712 16546
rect 338776 3398 338804 42162
rect 339420 5778 339448 85478
rect 340708 6662 340736 87774
rect 341628 85542 341656 87774
rect 342548 85542 342576 87774
rect 340788 85536 340840 85542
rect 340788 85478 340840 85484
rect 341616 85536 341668 85542
rect 341616 85478 341668 85484
rect 342168 85536 342220 85542
rect 342168 85478 342220 85484
rect 342536 85536 342588 85542
rect 342536 85478 342588 85484
rect 343456 85536 343508 85542
rect 343456 85478 343508 85484
rect 340800 6730 340828 85478
rect 340880 74112 340932 74118
rect 340880 74054 340932 74060
rect 340788 6724 340840 6730
rect 340788 6666 340840 6672
rect 340696 6656 340748 6662
rect 340696 6598 340748 6604
rect 339408 5772 339460 5778
rect 339408 5714 339460 5720
rect 339868 5636 339920 5642
rect 339868 5578 339920 5584
rect 338764 3392 338816 3398
rect 338764 3334 338816 3340
rect 339880 480 339908 5578
rect 340892 2038 340920 74054
rect 342180 5642 342208 85478
rect 343364 5840 343416 5846
rect 343364 5782 343416 5788
rect 342168 5636 342220 5642
rect 342168 5578 342220 5584
rect 340972 3052 341024 3058
rect 340972 2994 341024 3000
rect 340880 2032 340932 2038
rect 340880 1974 340932 1980
rect 340984 480 341012 2994
rect 342168 2032 342220 2038
rect 342168 1974 342220 1980
rect 342180 480 342208 1974
rect 343376 480 343404 5782
rect 343468 5778 343496 85478
rect 343560 5846 343588 87774
rect 344388 85542 344416 87774
rect 345216 85542 345244 87774
rect 344376 85536 344428 85542
rect 344376 85478 344428 85484
rect 344928 85536 344980 85542
rect 344928 85478 344980 85484
rect 345204 85536 345256 85542
rect 345204 85478 345256 85484
rect 344836 79348 344888 79354
rect 344836 79290 344888 79296
rect 344284 45008 344336 45014
rect 344284 44950 344336 44956
rect 343548 5840 343600 5846
rect 343548 5782 343600 5788
rect 343456 5772 343508 5778
rect 343456 5714 343508 5720
rect 344296 3058 344324 44950
rect 344848 6914 344876 79290
rect 344572 6886 344876 6914
rect 344284 3052 344336 3058
rect 344284 2994 344336 3000
rect 344572 480 344600 6886
rect 344940 5914 344968 85478
rect 346136 84194 346164 87774
rect 347056 85542 347084 87774
rect 347976 85542 348004 87774
rect 348896 86954 348924 87774
rect 348896 86926 349108 86954
rect 346308 85536 346360 85542
rect 346308 85478 346360 85484
rect 347044 85536 347096 85542
rect 347044 85478 347096 85484
rect 347688 85536 347740 85542
rect 347688 85478 347740 85484
rect 347964 85536 348016 85542
rect 347964 85478 348016 85484
rect 348976 85536 349028 85542
rect 348976 85478 349028 85484
rect 346136 84166 346256 84194
rect 346228 6866 346256 84166
rect 345756 6860 345808 6866
rect 345756 6802 345808 6808
rect 346216 6860 346268 6866
rect 346216 6802 346268 6808
rect 344928 5908 344980 5914
rect 344928 5850 344980 5856
rect 345768 480 345796 6802
rect 346320 6118 346348 85478
rect 347700 6798 347728 85478
rect 347688 6792 347740 6798
rect 347688 6734 347740 6740
rect 348988 6730 349016 85478
rect 348976 6724 349028 6730
rect 348976 6666 349028 6672
rect 349080 6662 349108 86926
rect 349816 85542 349844 87774
rect 350736 85542 350764 87774
rect 349804 85536 349856 85542
rect 349804 85478 349856 85484
rect 350448 85536 350500 85542
rect 350448 85478 350500 85484
rect 350724 85536 350776 85542
rect 350724 85478 350776 85484
rect 349804 65612 349856 65618
rect 349804 65554 349856 65560
rect 348792 6656 348844 6662
rect 348790 6624 348792 6633
rect 349068 6656 349120 6662
rect 348844 6624 348846 6633
rect 349068 6598 349120 6604
rect 348790 6559 348846 6568
rect 349252 6452 349304 6458
rect 349252 6394 349304 6400
rect 346308 6112 346360 6118
rect 346308 6054 346360 6060
rect 346952 5704 347004 5710
rect 346952 5646 347004 5652
rect 346964 480 346992 5646
rect 348056 3392 348108 3398
rect 348056 3334 348108 3340
rect 348068 480 348096 3334
rect 349264 480 349292 6394
rect 349816 3398 349844 65554
rect 350460 6458 350488 85478
rect 351656 85338 351684 87774
rect 351828 85536 351880 85542
rect 351828 85478 351880 85484
rect 351644 85332 351696 85338
rect 351644 85274 351696 85280
rect 350356 6452 350408 6458
rect 350356 6394 350408 6400
rect 350448 6452 350500 6458
rect 350448 6394 350500 6400
rect 349804 3392 349856 3398
rect 349804 3334 349856 3340
rect 350368 3346 350396 6394
rect 351840 6390 351868 85478
rect 352484 85066 352512 87774
rect 353404 85542 353432 87774
rect 353392 85536 353444 85542
rect 353392 85478 353444 85484
rect 354496 85536 354548 85542
rect 354496 85478 354548 85484
rect 352656 85332 352708 85338
rect 352656 85274 352708 85280
rect 352472 85060 352524 85066
rect 352472 85002 352524 85008
rect 352564 78056 352616 78062
rect 352564 77998 352616 78004
rect 351828 6384 351880 6390
rect 351828 6326 351880 6332
rect 352576 3398 352604 77998
rect 352668 17338 352696 85274
rect 352656 17332 352708 17338
rect 352656 17274 352708 17280
rect 354508 8974 354536 85478
rect 354496 8968 354548 8974
rect 354496 8910 354548 8916
rect 354600 8362 354628 87910
rect 355232 87802 355260 88049
rect 356152 87802 356180 88049
rect 357072 87802 357100 88049
rect 357992 87802 358020 88049
rect 358912 87802 358940 88049
rect 359740 87802 359768 88049
rect 360660 87802 360688 88049
rect 361580 87802 361608 88049
rect 362500 87802 362528 88049
rect 363420 87802 363448 88049
rect 364340 87802 364368 88049
rect 365260 87802 365288 88049
rect 366180 87802 366208 88049
rect 367008 87802 367036 88049
rect 355232 87774 355272 87802
rect 356152 87774 356192 87802
rect 357072 87774 357112 87802
rect 357992 87774 358032 87802
rect 358912 87774 358952 87802
rect 359740 87774 359780 87802
rect 360660 87774 360700 87802
rect 361580 87774 361620 87802
rect 362500 87774 362540 87802
rect 363420 87774 363460 87802
rect 364340 87774 364380 87802
rect 365260 87774 365300 87802
rect 366180 87774 366220 87802
rect 355244 85542 355272 87774
rect 356164 85542 356192 87774
rect 357084 87394 357112 87774
rect 357084 87366 357388 87394
rect 355232 85536 355284 85542
rect 355232 85478 355284 85484
rect 355968 85536 356020 85542
rect 355968 85478 356020 85484
rect 356152 85536 356204 85542
rect 356152 85478 356204 85484
rect 357256 85536 357308 85542
rect 357256 85478 357308 85484
rect 355980 8430 356008 85478
rect 357268 8498 357296 85478
rect 357360 8566 357388 87366
rect 358004 85542 358032 87774
rect 358924 85542 358952 87774
rect 359752 87394 359780 87774
rect 359752 87366 360148 87394
rect 357992 85536 358044 85542
rect 357992 85478 358044 85484
rect 358728 85536 358780 85542
rect 358728 85478 358780 85484
rect 358912 85536 358964 85542
rect 358912 85478 358964 85484
rect 360016 85536 360068 85542
rect 360016 85478 360068 85484
rect 358084 64320 358136 64326
rect 358084 64262 358136 64268
rect 357348 8560 357400 8566
rect 357348 8502 357400 8508
rect 357256 8492 357308 8498
rect 357256 8434 357308 8440
rect 355968 8424 356020 8430
rect 355968 8366 356020 8372
rect 354588 8356 354640 8362
rect 354588 8298 354640 8304
rect 354034 6624 354090 6633
rect 354034 6559 354090 6568
rect 352840 6316 352892 6322
rect 352840 6258 352892 6264
rect 351644 3392 351696 3398
rect 350368 3318 350488 3346
rect 351644 3334 351696 3340
rect 352564 3392 352616 3398
rect 352564 3334 352616 3340
rect 350460 480 350488 3318
rect 351656 480 351684 3334
rect 352852 480 352880 6258
rect 354048 480 354076 6559
rect 357532 5704 357584 5710
rect 357532 5646 357584 5652
rect 356336 5636 356388 5642
rect 356336 5578 356388 5584
rect 355232 3052 355284 3058
rect 355232 2994 355284 3000
rect 355244 480 355272 2994
rect 356348 480 356376 5578
rect 357544 480 357572 5646
rect 358096 3058 358124 64262
rect 358740 8634 358768 85478
rect 360028 8838 360056 85478
rect 360120 8906 360148 87366
rect 360672 85542 360700 87774
rect 361592 85542 361620 87774
rect 360660 85536 360712 85542
rect 360660 85478 360712 85484
rect 361488 85536 361540 85542
rect 361488 85478 361540 85484
rect 361580 85536 361632 85542
rect 361580 85478 361632 85484
rect 361500 9654 361528 85478
rect 362512 84194 362540 87774
rect 363432 85542 363460 87774
rect 364352 85542 364380 87774
rect 365272 86954 365300 87774
rect 365272 86926 365668 86954
rect 362868 85536 362920 85542
rect 362868 85478 362920 85484
rect 363420 85536 363472 85542
rect 363420 85478 363472 85484
rect 364248 85536 364300 85542
rect 364248 85478 364300 85484
rect 364340 85536 364392 85542
rect 364340 85478 364392 85484
rect 365536 85536 365588 85542
rect 365536 85478 365588 85484
rect 362512 84166 362816 84194
rect 361488 9648 361540 9654
rect 361488 9590 361540 9596
rect 362788 9518 362816 84166
rect 362880 9586 362908 85478
rect 362868 9580 362920 9586
rect 362868 9522 362920 9528
rect 362776 9512 362828 9518
rect 362776 9454 362828 9460
rect 364260 9450 364288 85478
rect 364248 9444 364300 9450
rect 364248 9386 364300 9392
rect 365548 9382 365576 85478
rect 365536 9376 365588 9382
rect 365536 9318 365588 9324
rect 365640 9110 365668 86926
rect 366192 85542 366220 87774
rect 366928 87774 367036 87802
rect 367928 87802 367956 88049
rect 368848 87802 368876 88049
rect 369768 87802 369796 88049
rect 367928 87774 367968 87802
rect 368848 87774 368888 87802
rect 366180 85536 366232 85542
rect 366180 85478 366232 85484
rect 365720 32496 365772 32502
rect 365720 32438 365772 32444
rect 365628 9104 365680 9110
rect 365628 9046 365680 9052
rect 360108 8900 360160 8906
rect 360108 8842 360160 8848
rect 360016 8832 360068 8838
rect 360016 8774 360068 8780
rect 358728 8628 358780 8634
rect 358728 8570 358780 8576
rect 359924 6248 359976 6254
rect 359924 6190 359976 6196
rect 358728 3732 358780 3738
rect 358728 3674 358780 3680
rect 358084 3052 358136 3058
rect 358084 2994 358136 3000
rect 358740 480 358768 3674
rect 359936 480 359964 6190
rect 363512 6180 363564 6186
rect 363512 6122 363564 6128
rect 361120 5772 361172 5778
rect 361120 5714 361172 5720
rect 361132 480 361160 5714
rect 362314 3360 362370 3369
rect 362314 3295 362370 3304
rect 362328 480 362356 3295
rect 363524 480 363552 6122
rect 364616 5840 364668 5846
rect 364616 5782 364668 5788
rect 364628 480 364656 5782
rect 365732 3398 365760 32438
rect 366928 9178 366956 87774
rect 367940 85542 367968 87774
rect 368860 85542 368888 87774
rect 369688 87774 369796 87802
rect 370688 87802 370716 88049
rect 371608 87802 371636 88049
rect 372528 87802 372556 88049
rect 373448 87802 373476 88049
rect 374276 87802 374304 88049
rect 375196 87802 375224 88049
rect 376116 87802 376144 88049
rect 377036 87802 377064 88049
rect 377956 87802 377984 88049
rect 378876 87802 378904 88049
rect 379796 87802 379824 88049
rect 380716 87802 380744 88049
rect 381636 87802 381664 88049
rect 382464 87802 382492 88049
rect 383384 87802 383412 88049
rect 384304 87802 384332 88049
rect 385224 87802 385252 88049
rect 386144 87938 386172 88049
rect 386144 87910 386368 87938
rect 370688 87774 370728 87802
rect 371608 87774 371648 87802
rect 372528 87774 372568 87802
rect 373448 87774 373488 87802
rect 374276 87774 374316 87802
rect 375196 87774 375328 87802
rect 376116 87774 376156 87802
rect 377036 87774 377076 87802
rect 377956 87774 377996 87802
rect 378876 87774 378916 87802
rect 379796 87774 379836 87802
rect 380716 87774 380756 87802
rect 381636 87774 381676 87802
rect 382464 87774 382504 87802
rect 383384 87774 383608 87802
rect 384304 87774 384344 87802
rect 385224 87774 385264 87802
rect 367008 85536 367060 85542
rect 367008 85478 367060 85484
rect 367928 85536 367980 85542
rect 367928 85478 367980 85484
rect 368388 85536 368440 85542
rect 368388 85478 368440 85484
rect 368848 85536 368900 85542
rect 368848 85478 368900 85484
rect 366916 9172 366968 9178
rect 366916 9114 366968 9120
rect 367020 7410 367048 85478
rect 368400 9042 368428 85478
rect 369688 10130 369716 87774
rect 370700 85542 370728 87774
rect 371620 85542 371648 87774
rect 369768 85536 369820 85542
rect 369768 85478 369820 85484
rect 370688 85536 370740 85542
rect 370688 85478 370740 85484
rect 371148 85536 371200 85542
rect 371148 85478 371200 85484
rect 371608 85536 371660 85542
rect 371608 85478 371660 85484
rect 372436 85536 372488 85542
rect 372436 85478 372488 85484
rect 369676 10124 369728 10130
rect 369676 10066 369728 10072
rect 369674 9208 369730 9217
rect 369674 9143 369730 9152
rect 369688 9110 369716 9143
rect 369780 9110 369808 85478
rect 369860 38004 369912 38010
rect 369860 37946 369912 37952
rect 369872 16574 369900 37946
rect 369872 16546 370636 16574
rect 369676 9104 369728 9110
rect 369676 9046 369728 9052
rect 369768 9104 369820 9110
rect 369768 9046 369820 9052
rect 368388 9036 368440 9042
rect 368388 8978 368440 8984
rect 367008 7404 367060 7410
rect 367008 7346 367060 7352
rect 368204 5908 368256 5914
rect 368204 5850 368256 5856
rect 365810 3496 365866 3505
rect 365810 3431 365866 3440
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 3431
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 368216 480 368244 5850
rect 369398 3632 369454 3641
rect 369398 3567 369454 3576
rect 369412 480 369440 3567
rect 370608 480 370636 16546
rect 371160 6934 371188 85478
rect 372448 10198 372476 85478
rect 372540 10266 372568 87774
rect 373460 84658 373488 87774
rect 374288 85542 374316 87774
rect 374276 85536 374328 85542
rect 374276 85478 374328 85484
rect 375196 85536 375248 85542
rect 375196 85478 375248 85484
rect 373448 84652 373500 84658
rect 373448 84594 373500 84600
rect 375208 73914 375236 85478
rect 375196 73908 375248 73914
rect 375196 73850 375248 73856
rect 375300 42158 375328 87774
rect 376128 85542 376156 87774
rect 377048 85542 377076 87774
rect 376116 85536 376168 85542
rect 376116 85478 376168 85484
rect 376668 85536 376720 85542
rect 376668 85478 376720 85484
rect 377036 85536 377088 85542
rect 377036 85478 377088 85484
rect 376024 84652 376076 84658
rect 376024 84594 376076 84600
rect 375288 42152 375340 42158
rect 375288 42094 375340 42100
rect 376036 39370 376064 84594
rect 376680 44946 376708 85478
rect 377968 50454 377996 87774
rect 378888 85542 378916 87774
rect 379808 85542 379836 87774
rect 378048 85536 378100 85542
rect 378048 85478 378100 85484
rect 378876 85536 378928 85542
rect 378876 85478 378928 85484
rect 379428 85536 379480 85542
rect 379428 85478 379480 85484
rect 379796 85536 379848 85542
rect 379796 85478 379848 85484
rect 377956 50448 378008 50454
rect 377956 50390 378008 50396
rect 378060 47666 378088 85478
rect 378048 47660 378100 47666
rect 378048 47602 378100 47608
rect 376668 44940 376720 44946
rect 376668 44882 376720 44888
rect 376760 42084 376812 42090
rect 376760 42026 376812 42032
rect 374000 39364 374052 39370
rect 374000 39306 374052 39312
rect 376024 39364 376076 39370
rect 376024 39306 376076 39312
rect 374012 16574 374040 39306
rect 376772 16574 376800 42026
rect 374012 16546 374132 16574
rect 376772 16546 377720 16574
rect 372528 10260 372580 10266
rect 372528 10202 372580 10208
rect 372436 10192 372488 10198
rect 372436 10134 372488 10140
rect 373906 9208 373962 9217
rect 373906 9143 373908 9152
rect 373960 9143 373962 9152
rect 373908 9114 373960 9120
rect 373724 9104 373776 9110
rect 373722 9072 373724 9081
rect 373776 9072 373778 9081
rect 373722 9007 373778 9016
rect 371148 6928 371200 6934
rect 371148 6870 371200 6876
rect 371700 6112 371752 6118
rect 371700 6054 371752 6060
rect 371712 480 371740 6054
rect 372894 3768 372950 3777
rect 372894 3703 372950 3712
rect 372908 480 372936 3703
rect 374104 480 374132 16546
rect 375288 6860 375340 6866
rect 375288 6802 375340 6808
rect 375300 480 375328 6802
rect 376484 3936 376536 3942
rect 376484 3878 376536 3884
rect 376496 480 376524 3878
rect 377692 480 377720 16546
rect 378876 6792 378928 6798
rect 378876 6734 378928 6740
rect 378888 480 378916 6734
rect 379440 6186 379468 85478
rect 379428 6180 379480 6186
rect 379428 6122 379480 6128
rect 380728 5642 380756 87774
rect 381648 85542 381676 87774
rect 382476 85542 382504 87774
rect 380808 85536 380860 85542
rect 380808 85478 380860 85484
rect 381636 85536 381688 85542
rect 381636 85478 381688 85484
rect 382188 85536 382240 85542
rect 382188 85478 382240 85484
rect 382464 85536 382516 85542
rect 382464 85478 382516 85484
rect 383476 85536 383528 85542
rect 383476 85478 383528 85484
rect 380820 6254 380848 85478
rect 380900 44872 380952 44878
rect 380900 44814 380952 44820
rect 380912 16574 380940 44814
rect 380912 16546 381216 16574
rect 380808 6248 380860 6254
rect 380808 6190 380860 6196
rect 380716 5636 380768 5642
rect 380716 5578 380768 5584
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379992 480 380020 3946
rect 381188 480 381216 16546
rect 382200 5710 382228 85478
rect 382372 6724 382424 6730
rect 382372 6666 382424 6672
rect 382188 5704 382240 5710
rect 382188 5646 382240 5652
rect 382384 480 382412 6666
rect 383488 5778 383516 85478
rect 383580 5846 383608 87774
rect 384316 85542 384344 87774
rect 385236 85542 385264 87774
rect 384304 85536 384356 85542
rect 384304 85478 384356 85484
rect 384948 85536 385000 85542
rect 384948 85478 385000 85484
rect 385224 85536 385276 85542
rect 385224 85478 385276 85484
rect 386236 85536 386288 85542
rect 386236 85478 386288 85484
rect 383660 47592 383712 47598
rect 383660 47534 383712 47540
rect 383672 16574 383700 47534
rect 383672 16546 384804 16574
rect 383568 5840 383620 5846
rect 383568 5782 383620 5788
rect 383476 5772 383528 5778
rect 383476 5714 383528 5720
rect 383660 5568 383712 5574
rect 383660 5510 383712 5516
rect 383672 5001 383700 5510
rect 383658 4992 383714 5001
rect 383658 4927 383714 4936
rect 383658 4856 383714 4865
rect 383658 4791 383714 4800
rect 383672 4146 383700 4791
rect 383660 4140 383712 4146
rect 383660 4082 383712 4088
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 383580 480 383608 4014
rect 384776 480 384804 16546
rect 384960 5914 384988 85478
rect 386248 16574 386276 85478
rect 386156 16546 386276 16574
rect 385960 6656 386012 6662
rect 385960 6598 386012 6604
rect 384948 5908 385000 5914
rect 384948 5850 385000 5856
rect 385972 480 386000 6598
rect 386156 6118 386184 16546
rect 386340 11778 386368 87910
rect 387064 87802 387092 88049
rect 387984 87802 388012 88049
rect 388904 87802 388932 88049
rect 389732 87802 389760 88049
rect 390652 87802 390680 88049
rect 391572 87802 391600 88049
rect 392492 87802 392520 88049
rect 393412 87802 393440 88049
rect 394332 87802 394360 88049
rect 395252 87802 395280 88049
rect 396172 87802 396200 88049
rect 397000 87802 397028 88049
rect 397920 87802 397948 88049
rect 398840 87802 398868 88049
rect 399760 87802 399788 88049
rect 400680 87802 400708 88049
rect 387064 87774 387104 87802
rect 387984 87774 388024 87802
rect 388904 87774 388944 87802
rect 389732 87774 389772 87802
rect 390652 87774 390692 87802
rect 391572 87774 391612 87802
rect 392492 87774 392532 87802
rect 393412 87774 393452 87802
rect 394332 87774 394372 87802
rect 395252 87774 395292 87802
rect 396172 87774 396212 87802
rect 397000 87774 397040 87802
rect 397920 87774 397960 87802
rect 398840 87774 398880 87802
rect 387076 85542 387104 87774
rect 387996 85542 388024 87774
rect 387064 85536 387116 85542
rect 387064 85478 387116 85484
rect 387708 85536 387760 85542
rect 387708 85478 387760 85484
rect 387984 85536 388036 85542
rect 387984 85478 388036 85484
rect 386248 11750 386368 11778
rect 386248 6866 386276 11750
rect 386236 6860 386288 6866
rect 386236 6802 386288 6808
rect 387720 6322 387748 85478
rect 388916 84194 388944 87774
rect 389744 85542 389772 87774
rect 390664 85542 390692 87774
rect 389088 85536 389140 85542
rect 389088 85478 389140 85484
rect 389732 85536 389784 85542
rect 389732 85478 389784 85484
rect 390468 85536 390520 85542
rect 390468 85478 390520 85484
rect 390652 85536 390704 85542
rect 390652 85478 390704 85484
rect 388916 84166 389036 84194
rect 387800 50380 387852 50386
rect 387800 50322 387852 50328
rect 387812 16574 387840 50322
rect 387812 16546 388300 16574
rect 387708 6316 387760 6322
rect 387708 6258 387760 6264
rect 386144 6112 386196 6118
rect 386144 6054 386196 6060
rect 387156 4140 387208 4146
rect 387156 4082 387208 4088
rect 387168 480 387196 4082
rect 388272 480 388300 16546
rect 389008 6798 389036 84166
rect 388996 6792 389048 6798
rect 388996 6734 389048 6740
rect 389100 6730 389128 85478
rect 389088 6724 389140 6730
rect 389088 6666 389140 6672
rect 390480 6662 390508 85478
rect 391584 84194 391612 87774
rect 392504 85542 392532 87774
rect 393424 85542 393452 87774
rect 391848 85536 391900 85542
rect 391848 85478 391900 85484
rect 392492 85536 392544 85542
rect 392492 85478 392544 85484
rect 393228 85536 393280 85542
rect 393228 85478 393280 85484
rect 393412 85536 393464 85542
rect 393412 85478 393464 85484
rect 391584 84166 391796 84194
rect 390560 14544 390612 14550
rect 390560 14486 390612 14492
rect 390468 6656 390520 6662
rect 390468 6598 390520 6604
rect 389456 6452 389508 6458
rect 389456 6394 389508 6400
rect 389468 480 389496 6394
rect 390572 3194 390600 14486
rect 391768 6458 391796 84166
rect 391756 6452 391808 6458
rect 391756 6394 391808 6400
rect 391860 6390 391888 85478
rect 391848 6384 391900 6390
rect 391848 6326 391900 6332
rect 393240 6322 393268 85478
rect 394344 84194 394372 87774
rect 395264 85542 395292 87774
rect 396184 85542 396212 87774
rect 397012 86170 397040 87774
rect 397012 86142 397408 86170
rect 394608 85536 394660 85542
rect 394608 85478 394660 85484
rect 395252 85536 395304 85542
rect 395252 85478 395304 85484
rect 395988 85536 396040 85542
rect 395988 85478 396040 85484
rect 396172 85536 396224 85542
rect 396172 85478 396224 85484
rect 397276 85536 397328 85542
rect 397276 85478 397328 85484
rect 394344 84166 394556 84194
rect 393320 8968 393372 8974
rect 393412 8968 393464 8974
rect 393320 8910 393372 8916
rect 393410 8936 393412 8945
rect 393464 8936 393466 8945
rect 393332 8809 393360 8910
rect 393410 8871 393466 8880
rect 393318 8800 393374 8809
rect 393318 8735 393374 8744
rect 394528 7342 394556 84166
rect 394516 7336 394568 7342
rect 394516 7278 394568 7284
rect 394620 6746 394648 85478
rect 394700 53100 394752 53106
rect 394700 53042 394752 53048
rect 394712 16574 394740 53042
rect 394712 16546 395384 16574
rect 394528 6718 394648 6746
rect 393044 6316 393096 6322
rect 393044 6258 393096 6264
rect 393228 6316 393280 6322
rect 393228 6258 393280 6264
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 390560 3188 390612 3194
rect 390560 3130 390612 3136
rect 390664 480 390692 3334
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 391860 480 391888 3130
rect 393056 480 393084 6258
rect 394528 6225 394556 6718
rect 394608 6656 394660 6662
rect 394608 6598 394660 6604
rect 394620 6254 394648 6598
rect 394608 6248 394660 6254
rect 394514 6216 394570 6225
rect 394608 6190 394660 6196
rect 394514 6151 394570 6160
rect 394240 3188 394292 3194
rect 394240 3130 394292 3136
rect 394252 480 394280 3130
rect 395356 480 395384 16546
rect 396000 7002 396028 85478
rect 396080 17332 396132 17338
rect 396080 17274 396132 17280
rect 396092 16574 396120 17274
rect 396092 16546 396580 16574
rect 395988 6996 396040 7002
rect 395988 6938 396040 6944
rect 396552 480 396580 16546
rect 397288 7206 397316 85478
rect 397380 7274 397408 86142
rect 397932 85542 397960 87774
rect 397920 85536 397972 85542
rect 397920 85478 397972 85484
rect 398748 85536 398800 85542
rect 398748 85478 398800 85484
rect 398104 85060 398156 85066
rect 398104 85002 398156 85008
rect 398116 13462 398144 85002
rect 398104 13456 398156 13462
rect 398104 13398 398156 13404
rect 398760 7342 398788 85478
rect 398852 10470 398880 87774
rect 399680 87774 399788 87802
rect 400600 87774 400708 87802
rect 401600 87802 401628 88049
rect 402520 87802 402548 88049
rect 402980 87848 403032 87854
rect 401600 87774 401640 87802
rect 402520 87774 402560 87802
rect 403440 87802 403468 88049
rect 404268 87854 404296 88049
rect 402980 87790 403032 87796
rect 399680 84194 399708 87774
rect 400600 84194 400628 87774
rect 401508 85536 401560 85542
rect 401508 85478 401560 85484
rect 398944 84166 399708 84194
rect 400232 84166 400628 84194
rect 398944 11762 398972 84166
rect 399024 55888 399076 55894
rect 399024 55830 399076 55836
rect 398932 11756 398984 11762
rect 398932 11698 398984 11704
rect 398840 10464 398892 10470
rect 398840 10406 398892 10412
rect 398656 7336 398708 7342
rect 398656 7278 398708 7284
rect 398748 7336 398800 7342
rect 398748 7278 398800 7284
rect 397368 7268 397420 7274
rect 397368 7210 397420 7216
rect 397276 7200 397328 7206
rect 397276 7142 397328 7148
rect 398668 7041 398696 7278
rect 398838 7168 398894 7177
rect 398838 7103 398894 7112
rect 398654 7032 398710 7041
rect 398852 7002 398880 7103
rect 398930 7032 398986 7041
rect 398654 6967 398710 6976
rect 398840 6996 398892 7002
rect 398930 6967 398932 6976
rect 398840 6938 398892 6944
rect 398984 6967 398986 6976
rect 398932 6938 398984 6944
rect 397736 3120 397788 3126
rect 397736 3062 397788 3068
rect 397748 480 397776 3062
rect 399036 2774 399064 55830
rect 400128 13456 400180 13462
rect 400128 13398 400180 13404
rect 398944 2746 399064 2774
rect 398944 480 398972 2746
rect 400140 480 400168 13398
rect 400232 11830 400260 84166
rect 401520 80714 401548 85478
rect 401612 84998 401640 87774
rect 402532 85542 402560 87774
rect 402520 85536 402572 85542
rect 402520 85478 402572 85484
rect 401600 84992 401652 84998
rect 401600 84934 401652 84940
rect 401508 80708 401560 80714
rect 401508 80650 401560 80656
rect 401600 18692 401652 18698
rect 401600 18634 401652 18640
rect 401612 16574 401640 18634
rect 401612 16546 402560 16574
rect 400220 11824 400272 11830
rect 400220 11766 400272 11772
rect 401324 3052 401376 3058
rect 401324 2994 401376 3000
rect 401336 480 401364 2994
rect 402532 480 402560 16546
rect 402992 3466 403020 87790
rect 403360 87774 403468 87802
rect 404256 87848 404308 87854
rect 405188 87802 405216 88049
rect 404256 87790 404308 87796
rect 405108 87774 405216 87802
rect 405740 87848 405792 87854
rect 406108 87802 406136 88049
rect 407028 87854 407056 88049
rect 405740 87790 405792 87796
rect 403360 84194 403388 87774
rect 405108 84194 405136 87774
rect 403084 84166 403388 84194
rect 404372 84166 405136 84194
rect 403084 61402 403112 84166
rect 403072 61396 403124 61402
rect 403072 61338 403124 61344
rect 403622 8800 403678 8809
rect 403622 8735 403678 8744
rect 402980 3460 403032 3466
rect 402980 3402 403032 3408
rect 403636 480 403664 8735
rect 404372 3534 404400 84166
rect 405752 3670 405780 87790
rect 406028 87774 406136 87802
rect 407016 87848 407068 87854
rect 407948 87802 407976 88049
rect 407016 87790 407068 87796
rect 407868 87774 407976 87802
rect 408500 87848 408552 87854
rect 408868 87802 408896 88049
rect 409788 87854 409816 88049
rect 408500 87790 408552 87796
rect 406028 84194 406056 87774
rect 407868 84194 407896 87774
rect 405844 84166 406056 84194
rect 407132 84166 407896 84194
rect 405740 3664 405792 3670
rect 405740 3606 405792 3612
rect 405844 3602 405872 84166
rect 405924 57248 405976 57254
rect 405924 57190 405976 57196
rect 405936 16574 405964 57190
rect 405936 16546 406056 16574
rect 405832 3596 405884 3602
rect 405832 3538 405884 3544
rect 404360 3528 404412 3534
rect 404360 3470 404412 3476
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 404832 480 404860 3402
rect 406028 480 406056 16546
rect 407132 10538 407160 84166
rect 408512 10674 408540 87790
rect 408788 87774 408896 87802
rect 409776 87848 409828 87854
rect 410708 87802 410736 88049
rect 411536 87802 411564 88049
rect 412456 87802 412484 88049
rect 413376 87802 413404 88049
rect 414296 87802 414324 88049
rect 415216 87802 415244 88049
rect 416136 87802 416164 88049
rect 417056 87802 417084 88049
rect 417976 87802 418004 88049
rect 418804 87802 418832 88049
rect 419724 87802 419752 88049
rect 420644 87802 420672 88049
rect 421564 87802 421592 88049
rect 409776 87790 409828 87796
rect 410628 87774 410736 87802
rect 411456 87774 411564 87802
rect 412376 87774 412484 87802
rect 413296 87774 413404 87802
rect 414216 87774 414324 87802
rect 415136 87774 415244 87802
rect 416056 87774 416164 87802
rect 416976 87774 417084 87802
rect 417896 87774 418004 87802
rect 418724 87774 418832 87802
rect 419552 87774 419752 87802
rect 420564 87774 420672 87802
rect 421484 87774 421592 87802
rect 422300 87848 422352 87854
rect 422484 87802 422512 88049
rect 423404 87854 423432 88049
rect 422300 87790 422352 87796
rect 408788 84194 408816 87774
rect 410628 84194 410656 87774
rect 411456 87496 411484 87774
rect 408604 84166 408816 84194
rect 409892 84166 410656 84194
rect 411272 87468 411484 87496
rect 408500 10668 408552 10674
rect 408500 10610 408552 10616
rect 408604 10606 408632 84166
rect 409604 13184 409656 13190
rect 409604 13126 409656 13132
rect 408592 10600 408644 10606
rect 408592 10542 408644 10548
rect 407120 10532 407172 10538
rect 407120 10474 407172 10480
rect 407212 8356 407264 8362
rect 407212 8298 407264 8304
rect 407224 480 407252 8298
rect 408314 7440 408370 7449
rect 408314 7375 408370 7384
rect 408328 7206 408356 7375
rect 408316 7200 408368 7206
rect 408408 7200 408460 7206
rect 408316 7142 408368 7148
rect 408406 7168 408408 7177
rect 408460 7168 408462 7177
rect 408406 7103 408462 7112
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 409616 480 409644 13126
rect 409892 10742 409920 84166
rect 411272 10810 411300 87468
rect 412376 84194 412404 87774
rect 413296 84194 413324 87774
rect 414216 87122 414244 87774
rect 411364 84166 412404 84194
rect 412652 84166 413324 84194
rect 414032 87094 414244 87122
rect 411364 11014 411392 84166
rect 412652 11898 412680 84166
rect 412732 60036 412784 60042
rect 412732 59978 412784 59984
rect 412744 16574 412772 59978
rect 412744 16546 413140 16574
rect 412640 11892 412692 11898
rect 412640 11834 412692 11840
rect 411352 11008 411404 11014
rect 411352 10950 411404 10956
rect 411260 10804 411312 10810
rect 411260 10746 411312 10752
rect 409880 10736 409932 10742
rect 409880 10678 409932 10684
rect 410800 8424 410852 8430
rect 410800 8366 410852 8372
rect 410812 480 410840 8366
rect 412640 7472 412692 7478
rect 412732 7472 412784 7478
rect 412640 7414 412692 7420
rect 412730 7440 412732 7449
rect 412784 7440 412786 7449
rect 412652 7313 412680 7414
rect 412730 7375 412786 7384
rect 412638 7304 412694 7313
rect 412638 7239 412694 7248
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 413112 480 413140 16546
rect 414032 12102 414060 87094
rect 415136 84194 415164 87774
rect 416056 84194 416084 87774
rect 416976 87122 417004 87774
rect 416792 87094 417004 87122
rect 416688 84992 416740 84998
rect 416688 84934 416740 84940
rect 414124 84166 415164 84194
rect 415412 84166 416084 84194
rect 414124 12170 414152 84166
rect 415412 12238 415440 84166
rect 415492 62824 415544 62830
rect 415492 62766 415544 62772
rect 415400 12232 415452 12238
rect 415400 12174 415452 12180
rect 414112 12164 414164 12170
rect 414112 12106 414164 12112
rect 414020 12096 414072 12102
rect 414020 12038 414072 12044
rect 414296 8492 414348 8498
rect 414296 8434 414348 8440
rect 414308 480 414336 8434
rect 415504 3670 415532 62766
rect 416700 6914 416728 84934
rect 416792 12306 416820 87094
rect 417896 84194 417924 87774
rect 418724 84194 418752 87774
rect 416884 84166 417924 84194
rect 418172 84166 418752 84194
rect 416884 12374 416912 84166
rect 418172 12442 418200 84166
rect 418160 12436 418212 12442
rect 418160 12378 418212 12384
rect 416872 12368 416924 12374
rect 416872 12310 416924 12316
rect 416780 12300 416832 12306
rect 416780 12242 416832 12248
rect 419552 11694 419580 87774
rect 420564 84194 420592 87774
rect 421484 84194 421512 87774
rect 419644 84166 420592 84194
rect 420932 84166 421512 84194
rect 419540 11688 419592 11694
rect 419540 11630 419592 11636
rect 419644 11626 419672 84166
rect 419724 21480 419776 21486
rect 419724 21422 419776 21428
rect 419736 16574 419764 21422
rect 419736 16546 420224 16574
rect 419632 11620 419684 11626
rect 419632 11562 419684 11568
rect 417884 8560 417936 8566
rect 417884 8502 417936 8508
rect 416608 6886 416728 6914
rect 415492 3664 415544 3670
rect 415492 3606 415544 3612
rect 416608 2990 416636 6886
rect 416688 3664 416740 3670
rect 416688 3606 416740 3612
rect 415492 2984 415544 2990
rect 415492 2926 415544 2932
rect 416596 2984 416648 2990
rect 416596 2926 416648 2932
rect 415504 480 415532 2926
rect 416700 480 416728 3606
rect 417896 480 417924 8502
rect 418988 2984 419040 2990
rect 418988 2926 419040 2932
rect 419000 480 419028 2926
rect 420196 480 420224 16546
rect 420932 11558 420960 84166
rect 420920 11552 420972 11558
rect 420920 11494 420972 11500
rect 422312 11286 422340 87790
rect 422404 87774 422512 87802
rect 423392 87848 423444 87854
rect 424324 87802 424352 88049
rect 425244 87802 425272 88049
rect 426072 87802 426100 88049
rect 426992 87802 427020 88049
rect 427912 87802 427940 88049
rect 428832 87802 428860 88049
rect 429752 87802 429780 88049
rect 423392 87790 423444 87796
rect 424244 87774 424352 87802
rect 425072 87774 425272 87802
rect 425992 87774 426100 87802
rect 426912 87774 427020 87802
rect 427832 87774 427940 87802
rect 428752 87774 428860 87802
rect 429672 87774 429780 87802
rect 430580 87848 430632 87854
rect 430580 87790 430632 87796
rect 430672 87802 430700 88049
rect 431592 87854 431620 88049
rect 431580 87848 431632 87854
rect 422404 11354 422432 87774
rect 423588 85060 423640 85066
rect 423588 85002 423640 85008
rect 422392 11348 422444 11354
rect 422392 11290 422444 11296
rect 422300 11280 422352 11286
rect 422300 11222 422352 11228
rect 421380 8628 421432 8634
rect 421380 8570 421432 8576
rect 421392 480 421420 8570
rect 423600 3670 423628 85002
rect 424244 84194 424272 87774
rect 423692 84166 424272 84194
rect 423692 11218 423720 84166
rect 425072 43450 425100 87774
rect 425992 84194 426020 87774
rect 426912 84194 426940 87774
rect 425164 84166 426020 84194
rect 426452 84166 426940 84194
rect 425164 54534 425192 84166
rect 425152 54528 425204 54534
rect 425152 54470 425204 54476
rect 425060 43444 425112 43450
rect 425060 43386 425112 43392
rect 423680 11212 423732 11218
rect 423680 11154 423732 11160
rect 426452 11150 426480 84166
rect 427832 33862 427860 87774
rect 428752 84194 428780 87774
rect 429672 84194 429700 87774
rect 427924 84166 428780 84194
rect 429212 84166 429700 84194
rect 427924 36582 427952 84166
rect 429212 40730 429240 84166
rect 430592 46374 430620 87790
rect 430672 87774 430712 87802
rect 432512 87802 432540 88049
rect 431580 87790 431632 87796
rect 430684 67046 430712 87774
rect 432432 87774 432540 87802
rect 433340 87802 433368 88049
rect 434260 87802 434288 88049
rect 435180 87802 435208 88049
rect 433340 87774 433380 87802
rect 432432 84194 432460 87774
rect 431972 84166 432460 84194
rect 430672 67040 430724 67046
rect 430672 66982 430724 66988
rect 430580 46368 430632 46374
rect 430580 46310 430632 46316
rect 429200 40724 429252 40730
rect 429200 40666 429252 40672
rect 427912 36576 427964 36582
rect 427912 36518 427964 36524
rect 427820 33856 427872 33862
rect 427820 33798 427872 33804
rect 431972 24206 432000 84166
rect 433352 49094 433380 87774
rect 434180 87774 434288 87802
rect 435100 87774 435208 87802
rect 436100 87802 436128 88049
rect 437020 87802 437048 88049
rect 437940 87802 437968 88049
rect 436100 87774 436140 87802
rect 434180 84194 434208 87774
rect 435100 84194 435128 87774
rect 436112 85542 436140 87774
rect 436940 87774 437048 87802
rect 437860 87774 437968 87802
rect 438860 87802 438888 88049
rect 439780 87802 439808 88049
rect 440608 87802 440636 88049
rect 438860 87774 438992 87802
rect 439780 87774 439820 87802
rect 435364 85536 435416 85542
rect 435364 85478 435416 85484
rect 436100 85536 436152 85542
rect 436100 85478 436152 85484
rect 433444 84166 434208 84194
rect 434732 84166 435128 84194
rect 433444 51814 433472 84166
rect 433432 51808 433484 51814
rect 433432 51750 433484 51756
rect 433340 49088 433392 49094
rect 433340 49030 433392 49036
rect 431960 24200 432012 24206
rect 431960 24142 432012 24148
rect 426440 11144 426492 11150
rect 426440 11086 426492 11092
rect 434732 11082 434760 84166
rect 435376 73846 435404 85478
rect 436940 84194 436968 87774
rect 437388 85128 437440 85134
rect 437388 85070 437440 85076
rect 436204 84166 436968 84194
rect 435364 73840 435416 73846
rect 435364 73782 435416 73788
rect 436204 58682 436232 84166
rect 436192 58676 436244 58682
rect 436192 58618 436244 58624
rect 434720 11076 434772 11082
rect 434720 11018 434772 11024
rect 432052 9648 432104 9654
rect 432052 9590 432104 9596
rect 428464 8900 428516 8906
rect 428464 8842 428516 8848
rect 424968 8832 425020 8838
rect 424968 8774 425020 8780
rect 423770 7304 423826 7313
rect 423770 7239 423826 7248
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 423588 3664 423640 3670
rect 423588 3606 423640 3612
rect 422588 480 422616 3606
rect 423784 480 423812 7239
rect 424980 480 425008 8774
rect 427268 7540 427320 7546
rect 427268 7482 427320 7488
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 426176 480 426204 2926
rect 427280 480 427308 7482
rect 428476 480 428504 8842
rect 430856 8288 430908 8294
rect 430856 8230 430908 8236
rect 429660 2916 429712 2922
rect 429660 2858 429712 2864
rect 429672 480 429700 2858
rect 430868 480 430896 8230
rect 432064 480 432092 9590
rect 435548 9580 435600 9586
rect 435548 9522 435600 9528
rect 434444 8084 434496 8090
rect 434444 8026 434496 8032
rect 433248 2848 433300 2854
rect 433248 2790 433300 2796
rect 433260 480 433288 2790
rect 434456 480 434484 8026
rect 435560 480 435588 9522
rect 437400 2854 437428 85070
rect 437860 84194 437888 87774
rect 438860 86148 438912 86154
rect 438860 86090 438912 86096
rect 437492 84166 437888 84194
rect 437492 76566 437520 84166
rect 437480 76560 437532 76566
rect 437480 76502 437532 76508
rect 438872 35290 438900 86090
rect 438964 53174 438992 87774
rect 439792 86154 439820 87774
rect 440528 87774 440636 87802
rect 441528 87802 441556 88049
rect 442448 87938 442476 88049
rect 442184 87910 442476 87938
rect 441528 87774 441568 87802
rect 439780 86148 439832 86154
rect 439780 86090 439832 86096
rect 439504 85536 439556 85542
rect 439504 85478 439556 85484
rect 438952 53168 439004 53174
rect 438952 53110 439004 53116
rect 438860 35284 438912 35290
rect 438860 35226 438912 35232
rect 439516 26994 439544 85478
rect 440528 84194 440556 87774
rect 441540 85542 441568 87774
rect 441528 85536 441580 85542
rect 441528 85478 441580 85484
rect 442184 84194 442212 87910
rect 443092 87848 443144 87854
rect 443092 87790 443144 87796
rect 443368 87802 443396 88049
rect 444288 87854 444316 88049
rect 444276 87848 444328 87854
rect 442264 85536 442316 85542
rect 442264 85478 442316 85484
rect 440344 84166 440556 84194
rect 441632 84166 442212 84194
rect 440344 83570 440372 84166
rect 440332 83564 440384 83570
rect 440332 83506 440384 83512
rect 441632 55962 441660 84166
rect 441620 55956 441672 55962
rect 441620 55898 441672 55904
rect 439504 26988 439556 26994
rect 439504 26930 439556 26936
rect 442276 22778 442304 85478
rect 443104 57322 443132 87790
rect 443368 87774 443408 87802
rect 445208 87802 445236 88049
rect 446128 87802 446156 88049
rect 444276 87790 444328 87796
rect 443380 85542 443408 87774
rect 445128 87774 445236 87802
rect 446048 87774 446156 87802
rect 447048 87802 447076 88049
rect 447876 87802 447904 88049
rect 447048 87774 447088 87802
rect 443368 85536 443420 85542
rect 443368 85478 443420 85484
rect 444288 85196 444340 85202
rect 444288 85138 444340 85144
rect 443092 57316 443144 57322
rect 443092 57258 443144 57264
rect 442264 22772 442316 22778
rect 442264 22714 442316 22720
rect 439136 9512 439188 9518
rect 439136 9454 439188 9460
rect 437940 8016 437992 8022
rect 437940 7958 437992 7964
rect 436744 2848 436796 2854
rect 436744 2790 436796 2796
rect 437388 2848 437440 2854
rect 437388 2790 437440 2796
rect 436756 480 436784 2790
rect 437952 480 437980 7958
rect 439148 480 439176 9454
rect 442632 9444 442684 9450
rect 442632 9386 442684 9392
rect 441528 7948 441580 7954
rect 441528 7890 441580 7896
rect 440332 2644 440384 2650
rect 440332 2586 440384 2592
rect 440344 480 440372 2586
rect 441540 480 441568 7890
rect 441710 3904 441766 3913
rect 441710 3839 441766 3848
rect 441724 2650 441752 3839
rect 441712 2644 441764 2650
rect 441712 2586 441764 2592
rect 442644 480 442672 9386
rect 444300 6914 444328 85138
rect 445128 84194 445156 87774
rect 446048 86954 446076 87774
rect 444392 84166 445156 84194
rect 445772 86926 446076 86954
rect 444392 82278 444420 84166
rect 444380 82272 444432 82278
rect 444380 82214 444432 82220
rect 445772 25702 445800 86926
rect 447060 86154 447088 87774
rect 447796 87774 447904 87802
rect 448520 87848 448572 87854
rect 448796 87802 448824 88049
rect 449716 87854 449744 88049
rect 448520 87790 448572 87796
rect 445852 86148 445904 86154
rect 445852 86090 445904 86096
rect 447048 86148 447100 86154
rect 447048 86090 447100 86096
rect 445864 60110 445892 86090
rect 447796 84194 447824 87774
rect 447152 84166 447824 84194
rect 445852 60104 445904 60110
rect 445852 60046 445904 60052
rect 447152 28422 447180 84166
rect 448532 29714 448560 87790
rect 448716 87774 448824 87802
rect 449704 87848 449756 87854
rect 450636 87802 450664 88049
rect 451556 87802 451584 88049
rect 452476 87802 452504 88049
rect 453396 87802 453424 88049
rect 449704 87790 449756 87796
rect 450556 87774 450664 87802
rect 451292 87774 451584 87802
rect 452396 87774 452504 87802
rect 453316 87774 453424 87802
rect 454040 87848 454092 87854
rect 454316 87802 454344 88049
rect 455144 87854 455172 88049
rect 454040 87790 454092 87796
rect 448716 84194 448744 87774
rect 450556 84194 450584 87774
rect 451188 85264 451240 85270
rect 451188 85206 451240 85212
rect 448624 84166 448744 84194
rect 449912 84166 450584 84194
rect 448624 62898 448652 84166
rect 448612 62892 448664 62898
rect 448612 62834 448664 62840
rect 449912 31142 449940 84166
rect 449900 31136 449952 31142
rect 449900 31078 449952 31084
rect 448520 29708 448572 29714
rect 448520 29650 448572 29656
rect 447140 28416 447192 28422
rect 447140 28358 447192 28364
rect 445760 25696 445812 25702
rect 445760 25638 445812 25644
rect 446220 9376 446272 9382
rect 446220 9318 446272 9324
rect 445024 7880 445076 7886
rect 445024 7822 445076 7828
rect 443840 6886 444328 6914
rect 443840 480 443868 6886
rect 445036 480 445064 7822
rect 446232 480 446260 9318
rect 449808 9172 449860 9178
rect 449808 9114 449860 9120
rect 448612 7812 448664 7818
rect 448612 7754 448664 7760
rect 447416 2644 447468 2650
rect 447416 2586 447468 2592
rect 447428 480 447456 2586
rect 448624 480 448652 7754
rect 449820 480 449848 9114
rect 451200 6914 451228 85206
rect 451292 39438 451320 87774
rect 452396 84194 452424 87774
rect 453316 84194 453344 87774
rect 451384 84166 452424 84194
rect 452672 84166 453344 84194
rect 451384 42226 451412 84166
rect 452672 45014 452700 84166
rect 454052 65618 454080 87790
rect 454236 87774 454344 87802
rect 455132 87848 455184 87854
rect 456064 87802 456092 88049
rect 455132 87790 455184 87796
rect 455984 87774 456092 87802
rect 456800 87848 456852 87854
rect 456984 87802 457012 88049
rect 457904 87854 457932 88049
rect 456800 87790 456852 87796
rect 454236 84194 454264 87774
rect 455328 85332 455380 85338
rect 455328 85274 455380 85280
rect 454144 84166 454264 84194
rect 454144 79354 454172 84166
rect 454132 79348 454184 79354
rect 454132 79290 454184 79296
rect 454040 65612 454092 65618
rect 454040 65554 454092 65560
rect 452660 45008 452712 45014
rect 452660 44950 452712 44956
rect 451372 42220 451424 42226
rect 451372 42162 451424 42168
rect 451280 39432 451332 39438
rect 451280 39374 451332 39380
rect 452108 7744 452160 7750
rect 452108 7686 452160 7692
rect 450924 6886 451228 6914
rect 450924 480 450952 6886
rect 451278 4040 451334 4049
rect 451278 3975 451334 3984
rect 451292 3738 451320 3975
rect 451372 3936 451424 3942
rect 451370 3904 451372 3913
rect 451424 3904 451426 3913
rect 451370 3839 451426 3848
rect 451280 3732 451332 3738
rect 451280 3674 451332 3680
rect 452120 480 452148 7686
rect 453304 7404 453356 7410
rect 453304 7346 453356 7352
rect 453316 480 453344 7346
rect 454406 3904 454462 3913
rect 454406 3839 454462 3848
rect 454420 3738 454448 3839
rect 455340 3738 455368 85274
rect 455984 84194 456012 87774
rect 455432 84166 456012 84194
rect 455432 78062 455460 84166
rect 455420 78056 455472 78062
rect 455420 77998 455472 78004
rect 455696 15904 455748 15910
rect 455696 15846 455748 15852
rect 455512 3936 455564 3942
rect 455510 3904 455512 3913
rect 455564 3904 455566 3913
rect 455510 3839 455566 3848
rect 454408 3732 454460 3738
rect 454408 3674 454460 3680
rect 454500 3732 454552 3738
rect 454500 3674 454552 3680
rect 455328 3732 455380 3738
rect 455328 3674 455380 3680
rect 454512 480 454540 3674
rect 455708 480 455736 15846
rect 456812 4049 456840 87790
rect 456904 87774 457012 87802
rect 457892 87848 457944 87854
rect 458824 87802 458852 88049
rect 457892 87790 457944 87796
rect 458744 87774 458852 87802
rect 459652 87848 459704 87854
rect 459652 87790 459704 87796
rect 459744 87802 459772 88049
rect 460664 87854 460692 88049
rect 460652 87848 460704 87854
rect 456904 64326 456932 87774
rect 458744 84194 458772 87774
rect 458192 84166 458772 84194
rect 456892 64320 456944 64326
rect 456892 64262 456944 64268
rect 456892 9104 456944 9110
rect 456892 9046 456944 9052
rect 456798 4040 456854 4049
rect 456798 3975 456854 3984
rect 456904 480 456932 9046
rect 458086 3904 458142 3913
rect 458086 3839 458142 3848
rect 458100 480 458128 3839
rect 458192 3369 458220 84166
rect 458272 65544 458324 65550
rect 458272 65486 458324 65492
rect 458284 16574 458312 65486
rect 458284 16546 459232 16574
rect 458178 3360 458234 3369
rect 458178 3295 458234 3304
rect 459204 480 459232 16546
rect 459664 3641 459692 87790
rect 459744 87774 459784 87802
rect 461584 87802 461612 88049
rect 462412 87802 462440 88049
rect 463332 87802 463360 88049
rect 464252 87802 464280 88049
rect 460652 87790 460704 87796
rect 459650 3632 459706 3641
rect 459650 3567 459706 3576
rect 459756 3505 459784 87774
rect 461504 87774 461612 87802
rect 462332 87774 462440 87802
rect 463252 87774 463360 87802
rect 464172 87774 464280 87802
rect 465172 87802 465200 88049
rect 466092 87802 466120 88049
rect 467012 87802 467040 88049
rect 465172 87774 465212 87802
rect 461504 84194 461532 87774
rect 462228 85536 462280 85542
rect 462228 85478 462280 85484
rect 460952 84166 461532 84194
rect 460388 9036 460440 9042
rect 460388 8978 460440 8984
rect 459742 3496 459798 3505
rect 459742 3431 459798 3440
rect 460400 480 460428 8978
rect 460662 4176 460718 4185
rect 460662 4111 460718 4120
rect 460570 4040 460626 4049
rect 460570 3975 460572 3984
rect 460624 3975 460626 3984
rect 460572 3946 460624 3952
rect 460676 3942 460704 4111
rect 460848 4004 460900 4010
rect 460848 3946 460900 3952
rect 460664 3936 460716 3942
rect 460860 3913 460888 3946
rect 460664 3878 460716 3884
rect 460846 3904 460902 3913
rect 460846 3839 460902 3848
rect 460952 3777 460980 84166
rect 461216 4140 461268 4146
rect 461216 4082 461268 4088
rect 461124 4072 461176 4078
rect 461122 4040 461124 4049
rect 461176 4040 461178 4049
rect 461228 4026 461256 4082
rect 461228 3998 461348 4026
rect 461122 3975 461178 3984
rect 460938 3768 460994 3777
rect 460938 3703 460994 3712
rect 461320 3194 461348 3998
rect 462240 3466 462268 85478
rect 462332 4185 462360 87774
rect 463252 84194 463280 87774
rect 464172 84194 464200 87774
rect 462424 84166 463280 84194
rect 463712 84166 464200 84194
rect 462318 4176 462374 4185
rect 462318 4111 462374 4120
rect 462424 4078 462452 84166
rect 462504 19984 462556 19990
rect 462504 19926 462556 19932
rect 462516 16574 462544 19926
rect 462516 16546 462820 16574
rect 462412 4072 462464 4078
rect 462412 4014 462464 4020
rect 461584 3460 461636 3466
rect 461584 3402 461636 3408
rect 462228 3460 462280 3466
rect 462228 3402 462280 3408
rect 462320 3460 462372 3466
rect 462320 3402 462372 3408
rect 461308 3188 461360 3194
rect 461308 3130 461360 3136
rect 460848 3120 460900 3126
rect 460938 3088 460994 3097
rect 460900 3068 460938 3074
rect 460848 3062 460938 3068
rect 460860 3046 460938 3062
rect 460938 3023 460994 3032
rect 461596 480 461624 3402
rect 462332 3097 462360 3402
rect 462318 3088 462374 3097
rect 462318 3023 462374 3032
rect 462792 480 462820 16546
rect 463712 3398 463740 84166
rect 463976 8968 464028 8974
rect 463976 8910 464028 8916
rect 463884 6248 463936 6254
rect 463882 6216 463884 6225
rect 463936 6216 463938 6225
rect 463882 6151 463938 6160
rect 463700 3392 463752 3398
rect 463700 3334 463752 3340
rect 463988 480 464016 8910
rect 465184 3346 465212 87774
rect 466012 87774 466120 87802
rect 466932 87774 467040 87802
rect 467932 87802 467960 88049
rect 468852 87802 468880 88049
rect 469680 87802 469708 88049
rect 467932 87774 467972 87802
rect 466012 84194 466040 87774
rect 466368 84788 466420 84794
rect 466368 84730 466420 84736
rect 465368 84166 466040 84194
rect 465264 68332 465316 68338
rect 465264 68274 465316 68280
rect 465092 3318 465212 3346
rect 465092 3194 465120 3318
rect 465080 3188 465132 3194
rect 465080 3130 465132 3136
rect 465172 3188 465224 3194
rect 465172 3130 465224 3136
rect 465184 480 465212 3130
rect 465276 2938 465304 68274
rect 465368 3126 465396 84166
rect 466380 3194 466408 84730
rect 466932 84194 466960 87774
rect 466472 84166 466960 84194
rect 466368 3188 466420 3194
rect 466368 3130 466420 3136
rect 465356 3120 465408 3126
rect 465356 3062 465408 3068
rect 466472 3058 466500 84166
rect 467472 10124 467524 10130
rect 467472 10066 467524 10072
rect 466460 3052 466512 3058
rect 466460 2994 466512 3000
rect 465276 2910 466316 2938
rect 466288 480 466316 2910
rect 467484 480 467512 10066
rect 467944 3466 467972 87774
rect 468772 87774 468880 87802
rect 469600 87774 469708 87802
rect 470600 87802 470628 88049
rect 471520 87802 471548 88049
rect 470600 87774 470640 87802
rect 468772 84194 468800 87774
rect 469128 84720 469180 84726
rect 469128 84662 469180 84668
rect 468036 84166 468800 84194
rect 468036 4146 468064 84166
rect 468024 4140 468076 4146
rect 468024 4082 468076 4088
rect 469140 3466 469168 84662
rect 469600 84194 469628 87774
rect 469232 84166 469628 84194
rect 469232 4078 469260 84166
rect 469312 71052 469364 71058
rect 469312 70994 469364 71000
rect 469324 16574 469352 70994
rect 469324 16546 469904 16574
rect 469220 4072 469272 4078
rect 469220 4014 469272 4020
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 468668 3460 468720 3466
rect 468668 3402 468720 3408
rect 469128 3460 469180 3466
rect 469128 3402 469180 3408
rect 468680 480 468708 3402
rect 469876 480 469904 16546
rect 470612 3534 470640 87774
rect 471440 87774 471548 87802
rect 472440 87802 472468 88049
rect 473360 87802 473388 88049
rect 474280 87802 474308 88049
rect 475200 87802 475228 88049
rect 472440 87774 472480 87802
rect 473360 87774 473400 87802
rect 474280 87774 474320 87802
rect 471440 84194 471468 87774
rect 472452 84998 472480 87774
rect 472440 84992 472492 84998
rect 472440 84934 472492 84940
rect 473268 84992 473320 84998
rect 473268 84934 473320 84940
rect 470704 84166 471468 84194
rect 470704 16574 470732 84166
rect 470704 16546 470824 16574
rect 470690 4856 470746 4865
rect 470690 4791 470746 4800
rect 470704 4078 470732 4791
rect 470692 4072 470744 4078
rect 470692 4014 470744 4020
rect 470796 3602 470824 16546
rect 471060 7404 471112 7410
rect 471060 7346 471112 7352
rect 470784 3596 470836 3602
rect 470784 3538 470836 3544
rect 470600 3528 470652 3534
rect 470600 3470 470652 3476
rect 471072 480 471100 7346
rect 473280 3194 473308 84934
rect 473372 84194 473400 87774
rect 474292 85066 474320 87774
rect 475120 87774 475228 87802
rect 476120 87802 476148 88049
rect 476948 87802 476976 88049
rect 476120 87774 476160 87802
rect 474280 85060 474332 85066
rect 474280 85002 474332 85008
rect 475120 84194 475148 87774
rect 476028 85060 476080 85066
rect 476028 85002 476080 85008
rect 473372 84166 473584 84194
rect 473452 32428 473504 32434
rect 473452 32370 473504 32376
rect 472256 3188 472308 3194
rect 472256 3130 472308 3136
rect 473268 3188 473320 3194
rect 473268 3130 473320 3136
rect 472268 480 472296 3130
rect 473464 480 473492 32370
rect 473556 3670 473584 84166
rect 474844 84166 475148 84194
rect 474556 10192 474608 10198
rect 474556 10134 474608 10140
rect 473544 3664 473596 3670
rect 473544 3606 473596 3612
rect 474568 480 474596 10134
rect 474844 2990 474872 84166
rect 476040 6914 476068 85002
rect 475764 6886 476068 6914
rect 474832 2984 474884 2990
rect 474832 2926 474884 2932
rect 475764 480 475792 6886
rect 476132 2922 476160 87774
rect 476868 87774 476976 87802
rect 477868 87802 477896 88049
rect 478788 87802 478816 88049
rect 477868 87774 477908 87802
rect 476868 84194 476896 87774
rect 477880 85134 477908 87774
rect 478708 87774 478816 87802
rect 479708 87802 479736 88049
rect 480628 87802 480656 88049
rect 479708 87774 479748 87802
rect 477868 85128 477920 85134
rect 477868 85070 477920 85076
rect 478708 84194 478736 87774
rect 479720 85202 479748 87774
rect 480548 87774 480656 87802
rect 481548 87802 481576 88049
rect 482468 87802 482496 88049
rect 483388 87802 483416 88049
rect 481548 87774 481588 87802
rect 482468 87774 482508 87802
rect 479708 85196 479760 85202
rect 479708 85138 479760 85144
rect 480168 85128 480220 85134
rect 480168 85070 480220 85076
rect 476224 84166 476896 84194
rect 477696 84166 478736 84194
rect 476120 2916 476172 2922
rect 476120 2858 476172 2864
rect 476224 2854 476252 84166
rect 476304 37936 476356 37942
rect 476304 37878 476356 37884
rect 476316 16574 476344 37878
rect 476316 16546 476988 16574
rect 476212 2848 476264 2854
rect 476212 2790 476264 2796
rect 476960 480 476988 16546
rect 477592 10260 477644 10266
rect 477592 10202 477644 10208
rect 477604 3482 477632 10202
rect 477696 3738 477724 84166
rect 477684 3732 477736 3738
rect 477684 3674 477736 3680
rect 480180 3534 480208 85070
rect 480548 84194 480576 87774
rect 481560 85270 481588 87774
rect 482480 85338 482508 87774
rect 483308 87774 483416 87802
rect 484308 87802 484336 88049
rect 485136 87802 485164 88049
rect 486056 87802 486084 88049
rect 486976 87802 487004 88049
rect 487896 87802 487924 88049
rect 488816 87802 488844 88049
rect 489736 87802 489764 88049
rect 490656 87802 490684 88049
rect 491576 87802 491604 88049
rect 484308 87774 484348 87802
rect 485136 87774 485176 87802
rect 486056 87774 486096 87802
rect 486976 87774 487016 87802
rect 487896 87774 487936 87802
rect 488816 87774 488856 87802
rect 489736 87774 489776 87802
rect 490656 87774 490696 87802
rect 482468 85332 482520 85338
rect 482468 85274 482520 85280
rect 482928 85332 482980 85338
rect 482928 85274 482980 85280
rect 481548 85264 481600 85270
rect 481548 85206 481600 85212
rect 480456 84166 480576 84194
rect 480456 16574 480484 84166
rect 481640 39364 481692 39370
rect 481640 39306 481692 39312
rect 481652 16574 481680 39306
rect 480456 16546 480668 16574
rect 481652 16546 481772 16574
rect 480352 14476 480404 14482
rect 480352 14418 480404 14424
rect 480364 5114 480392 14418
rect 480364 5086 480576 5114
rect 480350 4992 480406 5001
rect 480350 4927 480406 4936
rect 480258 4856 480314 4865
rect 480364 4826 480392 4927
rect 480258 4791 480260 4800
rect 480312 4791 480314 4800
rect 480352 4820 480404 4826
rect 480260 4762 480312 4768
rect 480352 4762 480404 4768
rect 479340 3528 479392 3534
rect 477604 3454 478184 3482
rect 479340 3470 479392 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 478156 480 478184 3454
rect 479352 480 479380 3470
rect 480548 480 480576 5086
rect 480640 3942 480668 16546
rect 480628 3936 480680 3942
rect 480628 3878 480680 3884
rect 481744 480 481772 16546
rect 482940 6914 482968 85274
rect 483308 84194 483336 87774
rect 484320 85542 484348 87774
rect 484308 85536 484360 85542
rect 484308 85478 484360 85484
rect 485148 84794 485176 87774
rect 485136 84788 485188 84794
rect 485136 84730 485188 84736
rect 486068 84726 486096 87774
rect 486988 84998 487016 87774
rect 487908 85066 487936 87774
rect 488828 85134 488856 87774
rect 489748 85338 489776 87774
rect 489736 85332 489788 85338
rect 489736 85274 489788 85280
rect 488816 85128 488868 85134
rect 488816 85070 488868 85076
rect 487896 85060 487948 85066
rect 487896 85002 487948 85008
rect 486976 84992 487028 84998
rect 486976 84934 487028 84940
rect 486056 84720 486108 84726
rect 486056 84662 486108 84668
rect 490668 84250 490696 87774
rect 491496 87774 491604 87802
rect 492404 87802 492432 88049
rect 493324 87802 493352 88049
rect 494244 87802 494272 88049
rect 495164 87802 495192 88049
rect 496084 87802 496112 88049
rect 497004 87802 497032 88049
rect 497924 87802 497952 88049
rect 498844 87802 498872 88049
rect 499672 87802 499700 88049
rect 500592 87802 500620 88049
rect 501512 87802 501540 88049
rect 502432 87802 502460 88049
rect 503352 87802 503380 88049
rect 504272 87802 504300 88049
rect 505192 87802 505220 88049
rect 506112 87802 506140 88049
rect 506940 87802 506968 88049
rect 507860 87802 507888 88049
rect 508780 87802 508808 88049
rect 509700 87802 509728 88049
rect 510620 87802 510648 88049
rect 511540 87802 511568 88049
rect 512460 87802 512488 88049
rect 513380 87802 513408 88049
rect 514208 87802 514236 88049
rect 515128 87802 515156 88049
rect 516048 87802 516076 88049
rect 492404 87774 492444 87802
rect 493324 87774 493364 87802
rect 494244 87774 494284 87802
rect 495164 87774 495204 87802
rect 496084 87774 496124 87802
rect 497004 87774 497044 87802
rect 497924 87774 497964 87802
rect 498844 87774 498884 87802
rect 499672 87774 499712 87802
rect 500592 87774 500632 87802
rect 501512 87774 501552 87802
rect 502432 87774 502472 87802
rect 503352 87774 503392 87802
rect 504272 87774 504312 87802
rect 505192 87774 505232 87802
rect 506112 87774 506152 87802
rect 506940 87774 506980 87802
rect 507860 87774 507900 87802
rect 508780 87774 508820 87802
rect 509700 87774 509740 87802
rect 510620 87774 510660 87802
rect 511540 87774 511580 87802
rect 512460 87774 512500 87802
rect 513380 87774 513420 87802
rect 514208 87774 514248 87802
rect 515128 87774 515168 87802
rect 483216 84166 483336 84194
rect 487068 84244 487120 84250
rect 487068 84186 487120 84192
rect 490656 84244 490708 84250
rect 491496 84194 491524 87774
rect 490656 84186 490708 84192
rect 483112 83496 483164 83502
rect 483112 83438 483164 83444
rect 482848 6886 482968 6914
rect 482848 480 482876 6886
rect 483124 3482 483152 83438
rect 483216 4010 483244 84166
rect 484400 73908 484452 73914
rect 484400 73850 484452 73856
rect 484412 16574 484440 73850
rect 485044 50448 485096 50454
rect 485044 50390 485096 50396
rect 484412 16546 484992 16574
rect 483204 4004 483256 4010
rect 483204 3946 483256 3952
rect 484964 3482 484992 16546
rect 485056 3602 485084 50390
rect 485044 3596 485096 3602
rect 485044 3538 485096 3544
rect 487080 3534 487108 84186
rect 491220 84166 491524 84194
rect 492416 84194 492444 87774
rect 493336 85542 493364 87774
rect 494256 85542 494284 87774
rect 493324 85536 493376 85542
rect 493324 85478 493376 85484
rect 493968 85536 494020 85542
rect 493968 85478 494020 85484
rect 494244 85536 494296 85542
rect 494244 85478 494296 85484
rect 492416 84166 492812 84194
rect 487160 80776 487212 80782
rect 487160 80718 487212 80724
rect 487172 16574 487200 80718
rect 487804 47660 487856 47666
rect 487804 47602 487856 47608
rect 487172 16546 487660 16574
rect 486424 3528 486476 3534
rect 483124 3454 484072 3482
rect 484964 3454 485268 3482
rect 486424 3470 486476 3476
rect 487068 3528 487120 3534
rect 487068 3470 487120 3476
rect 484044 480 484072 3454
rect 485240 480 485268 3454
rect 486436 480 486464 3470
rect 487632 480 487660 16546
rect 487816 3534 487844 47602
rect 489184 44940 489236 44946
rect 489184 44882 489236 44888
rect 488540 42152 488592 42158
rect 488540 42094 488592 42100
rect 488552 16574 488580 42094
rect 488552 16546 488856 16574
rect 487804 3528 487856 3534
rect 487804 3470 487856 3476
rect 488828 480 488856 16546
rect 489196 4010 489224 44882
rect 489920 17264 489972 17270
rect 489920 17206 489972 17212
rect 489932 11762 489960 17206
rect 489920 11756 489972 11762
rect 489920 11698 489972 11704
rect 491116 11756 491168 11762
rect 491116 11698 491168 11704
rect 489918 5128 489974 5137
rect 489918 5063 489974 5072
rect 489826 4992 489882 5001
rect 489826 4927 489882 4936
rect 489840 4826 489868 4927
rect 489932 4826 489960 5063
rect 489828 4820 489880 4826
rect 489828 4762 489880 4768
rect 489920 4820 489972 4826
rect 489920 4762 489972 4768
rect 489184 4004 489236 4010
rect 489184 3946 489236 3952
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 489932 480 489960 3538
rect 491128 480 491156 11698
rect 491220 3602 491248 84166
rect 492784 16574 492812 84166
rect 492784 16546 493548 16574
rect 492312 4004 492364 4010
rect 492312 3946 492364 3952
rect 491208 3596 491260 3602
rect 491208 3538 491260 3544
rect 492324 480 492352 3946
rect 493520 480 493548 16546
rect 493980 3534 494008 85478
rect 495176 84998 495204 87774
rect 496096 85542 496124 87774
rect 497016 85542 497044 87774
rect 495348 85536 495400 85542
rect 495348 85478 495400 85484
rect 496084 85536 496136 85542
rect 496084 85478 496136 85484
rect 496728 85536 496780 85542
rect 496728 85478 496780 85484
rect 497004 85536 497056 85542
rect 497004 85478 497056 85484
rect 495164 84992 495216 84998
rect 495164 84934 495216 84940
rect 494060 18624 494112 18630
rect 494060 18566 494112 18572
rect 494072 16574 494100 18566
rect 494072 16546 494744 16574
rect 493968 3528 494020 3534
rect 493968 3470 494020 3476
rect 494716 480 494744 16546
rect 495360 3738 495388 85478
rect 496740 3942 496768 85478
rect 497936 84194 497964 87774
rect 498856 85542 498884 87774
rect 499684 85542 499712 87774
rect 500604 87258 500632 87774
rect 500604 87230 500908 87258
rect 498108 85536 498160 85542
rect 498108 85478 498160 85484
rect 498844 85536 498896 85542
rect 498844 85478 498896 85484
rect 499488 85536 499540 85542
rect 499488 85478 499540 85484
rect 499672 85536 499724 85542
rect 499672 85478 499724 85484
rect 500776 85536 500828 85542
rect 500776 85478 500828 85484
rect 497936 84166 498056 84194
rect 498028 4010 498056 84166
rect 498016 4004 498068 4010
rect 498016 3946 498068 3952
rect 496728 3936 496780 3942
rect 496728 3878 496780 3884
rect 495348 3732 495400 3738
rect 495348 3674 495400 3680
rect 498120 3670 498148 85478
rect 498292 21412 498344 21418
rect 498292 21354 498344 21360
rect 498304 6914 498332 21354
rect 499500 6914 499528 85478
rect 498212 6886 498332 6914
rect 499316 6886 499528 6914
rect 498108 3664 498160 3670
rect 498108 3606 498160 3612
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 495900 3460 495952 3466
rect 495900 3402 495952 3408
rect 495912 480 495940 3402
rect 497108 480 497136 3470
rect 498212 480 498240 6886
rect 499316 3602 499344 6886
rect 499672 5568 499724 5574
rect 499670 5536 499672 5545
rect 499764 5568 499816 5574
rect 499724 5536 499726 5545
rect 499764 5510 499816 5516
rect 499670 5471 499726 5480
rect 499776 5001 499804 5510
rect 499394 4992 499450 5001
rect 499394 4927 499450 4936
rect 499762 4992 499818 5001
rect 499762 4927 499818 4936
rect 499408 4826 499436 4927
rect 499486 4856 499542 4865
rect 499396 4820 499448 4826
rect 499486 4791 499488 4800
rect 499396 4762 499448 4768
rect 499540 4791 499542 4800
rect 499488 4762 499540 4768
rect 500592 3732 500644 3738
rect 500592 3674 500644 3680
rect 499304 3596 499356 3602
rect 499304 3538 499356 3544
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500604 480 500632 3674
rect 500788 3534 500816 85478
rect 500776 3528 500828 3534
rect 500776 3470 500828 3476
rect 500880 3466 500908 87230
rect 501524 85542 501552 87774
rect 502444 85542 502472 87774
rect 503364 87258 503392 87774
rect 503364 87230 503668 87258
rect 501512 85536 501564 85542
rect 501512 85478 501564 85484
rect 502248 85536 502300 85542
rect 502248 85478 502300 85484
rect 502432 85536 502484 85542
rect 502432 85478 502484 85484
rect 503536 85536 503588 85542
rect 503536 85478 503588 85484
rect 500960 24132 501012 24138
rect 500960 24074 501012 24080
rect 500972 16574 501000 24074
rect 500972 16546 501828 16574
rect 500868 3460 500920 3466
rect 500868 3402 500920 3408
rect 501800 480 501828 16546
rect 502260 6914 502288 85478
rect 502076 6886 502288 6914
rect 502076 2854 502104 6886
rect 502156 6180 502208 6186
rect 502156 6122 502208 6128
rect 502168 6066 502196 6122
rect 502168 6038 503024 6066
rect 502064 2848 502116 2854
rect 502064 2790 502116 2796
rect 502996 480 503024 6038
rect 503548 2922 503576 85478
rect 503640 2990 503668 87230
rect 504284 85542 504312 87774
rect 505204 85542 505232 87774
rect 506124 87258 506152 87774
rect 506124 87230 506428 87258
rect 504272 85536 504324 85542
rect 504272 85478 504324 85484
rect 505008 85536 505060 85542
rect 505008 85478 505060 85484
rect 505192 85536 505244 85542
rect 505192 85478 505244 85484
rect 506296 85536 506348 85542
rect 506296 85478 506348 85484
rect 503812 84992 503864 84998
rect 503812 84934 503864 84940
rect 503824 16574 503852 84934
rect 503824 16546 504220 16574
rect 503628 2984 503680 2990
rect 503628 2926 503680 2932
rect 503536 2916 503588 2922
rect 503536 2858 503588 2864
rect 504192 480 504220 16546
rect 505020 3058 505048 85478
rect 505100 26920 505152 26926
rect 505100 26862 505152 26868
rect 505112 16574 505140 26862
rect 505112 16546 505416 16574
rect 505008 3052 505060 3058
rect 505008 2994 505060 3000
rect 505388 480 505416 16546
rect 506308 3126 506336 85478
rect 506400 3194 506428 87230
rect 506952 85542 506980 87774
rect 507872 85542 507900 87774
rect 508792 87530 508820 87774
rect 508792 87502 509188 87530
rect 506940 85536 506992 85542
rect 506940 85478 506992 85484
rect 507768 85536 507820 85542
rect 507768 85478 507820 85484
rect 507860 85536 507912 85542
rect 507860 85478 507912 85484
rect 509056 85536 509108 85542
rect 509056 85478 509108 85484
rect 506478 5536 506534 5545
rect 506478 5471 506534 5480
rect 506388 3188 506440 3194
rect 506388 3130 506440 3136
rect 506296 3120 506348 3126
rect 506296 3062 506348 3068
rect 506492 480 506520 5471
rect 507676 3936 507728 3942
rect 507676 3878 507728 3884
rect 507688 480 507716 3878
rect 507780 3398 507808 85478
rect 507860 29640 507912 29646
rect 507860 29582 507912 29588
rect 507872 16574 507900 29582
rect 507872 16546 508912 16574
rect 507768 3392 507820 3398
rect 507768 3334 507820 3340
rect 508884 480 508912 16546
rect 509068 3942 509096 85478
rect 509160 4078 509188 87502
rect 509712 85542 509740 87774
rect 510632 85542 510660 87774
rect 511552 87394 511580 87774
rect 511552 87366 511948 87394
rect 509700 85536 509752 85542
rect 509700 85478 509752 85484
rect 510528 85536 510580 85542
rect 510528 85478 510580 85484
rect 510620 85536 510672 85542
rect 510620 85478 510672 85484
rect 511816 85536 511868 85542
rect 511816 85478 511868 85484
rect 510068 5636 510120 5642
rect 510068 5578 510120 5584
rect 509240 5024 509292 5030
rect 509238 4992 509240 5001
rect 509292 4992 509294 5001
rect 509238 4927 509294 4936
rect 509148 4072 509200 4078
rect 509148 4014 509200 4020
rect 509056 3936 509108 3942
rect 509056 3878 509108 3884
rect 510080 480 510108 5578
rect 510540 4146 510568 85478
rect 510528 4140 510580 4146
rect 510528 4082 510580 4088
rect 511828 3738 511856 85478
rect 511920 3913 511948 87366
rect 512472 85542 512500 87774
rect 512460 85536 512512 85542
rect 512460 85478 512512 85484
rect 513288 85536 513340 85542
rect 513288 85478 513340 85484
rect 512458 4992 512514 5001
rect 512458 4927 512514 4936
rect 511906 3904 511962 3913
rect 511906 3839 511962 3848
rect 511264 3732 511316 3738
rect 511264 3674 511316 3680
rect 511816 3732 511868 3738
rect 511816 3674 511868 3680
rect 511276 480 511304 3674
rect 512472 480 512500 4927
rect 513300 3777 513328 85478
rect 513392 85338 513420 87774
rect 514220 85542 514248 87774
rect 515140 85542 515168 87774
rect 515968 87774 516076 87802
rect 516968 87802 516996 88049
rect 517888 87802 517916 88049
rect 516968 87774 517008 87802
rect 517888 87774 517928 87802
rect 514208 85536 514260 85542
rect 514208 85478 514260 85484
rect 514668 85536 514720 85542
rect 514668 85478 514720 85484
rect 515128 85536 515180 85542
rect 515128 85478 515180 85484
rect 513380 85332 513432 85338
rect 513380 85274 513432 85280
rect 514576 85332 514628 85338
rect 514576 85274 514628 85280
rect 513564 5704 513616 5710
rect 513564 5646 513616 5652
rect 513286 3768 513342 3777
rect 513286 3703 513342 3712
rect 513576 480 513604 5646
rect 514588 5574 514616 85274
rect 514576 5568 514628 5574
rect 514576 5510 514628 5516
rect 514680 3505 514708 85478
rect 515968 6914 515996 87774
rect 516980 85542 517008 87774
rect 517900 85542 517928 87774
rect 516048 85536 516100 85542
rect 516048 85478 516100 85484
rect 516968 85536 517020 85542
rect 516968 85478 517020 85484
rect 517428 85536 517480 85542
rect 517428 85478 517480 85484
rect 517888 85536 517940 85542
rect 517888 85478 517940 85484
rect 518808 85536 518860 85542
rect 518808 85478 518860 85484
rect 515876 6886 515996 6914
rect 514760 3664 514812 3670
rect 514760 3606 514812 3612
rect 514666 3496 514722 3505
rect 514666 3431 514722 3440
rect 514772 480 514800 3606
rect 515876 3369 515904 6886
rect 515956 4004 516008 4010
rect 515956 3946 516008 3952
rect 515862 3360 515918 3369
rect 515862 3295 515918 3304
rect 515968 480 515996 3946
rect 516060 3670 516088 85478
rect 517152 5772 517204 5778
rect 517152 5714 517204 5720
rect 516230 3768 516286 3777
rect 516230 3703 516232 3712
rect 516284 3703 516286 3712
rect 516232 3674 516284 3680
rect 516048 3664 516100 3670
rect 516048 3606 516100 3612
rect 517164 480 517192 5714
rect 517440 3641 517468 85478
rect 518622 3904 518678 3913
rect 518622 3839 518678 3848
rect 518636 3738 518664 3839
rect 518820 3777 518848 85478
rect 520936 5846 520964 88839
rect 521028 20602 521056 99311
rect 521120 33114 521148 110599
rect 521212 46918 521240 122023
rect 521304 60722 521332 133447
rect 521396 73166 521424 144735
rect 521488 86970 521516 156159
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113076 580224 113082
rect 580172 113018 580224 113024
rect 580184 112849 580212 113018
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100564 580224 100570
rect 580172 100506 580224 100512
rect 580184 99521 580212 100506
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 521476 86964 521528 86970
rect 521476 86906 521528 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 572720 77988 572772 77994
rect 572720 77930 572772 77936
rect 568580 75200 568632 75206
rect 568580 75142 568632 75148
rect 521384 73160 521436 73166
rect 521384 73102 521436 73108
rect 521292 60716 521344 60722
rect 521292 60658 521344 60664
rect 521200 46912 521252 46918
rect 521200 46854 521252 46860
rect 521108 33108 521160 33114
rect 521108 33050 521160 33056
rect 521016 20596 521068 20602
rect 521016 20538 521068 20544
rect 568592 16574 568620 75142
rect 568592 16546 569172 16574
rect 566832 7200 566884 7206
rect 566832 7142 566884 7148
rect 563244 6996 563296 7002
rect 563244 6938 563296 6944
rect 531320 6860 531372 6866
rect 531320 6802 531372 6808
rect 527824 6112 527876 6118
rect 527824 6054 527876 6060
rect 524236 5908 524288 5914
rect 524236 5850 524288 5856
rect 520740 5840 520792 5846
rect 520740 5782 520792 5788
rect 520924 5840 520976 5846
rect 520924 5782 520976 5788
rect 519544 4208 519596 4214
rect 519544 4150 519596 4156
rect 518806 3768 518862 3777
rect 518624 3732 518676 3738
rect 518806 3703 518862 3712
rect 518990 3768 519046 3777
rect 518990 3703 519046 3712
rect 518624 3674 518676 3680
rect 517426 3632 517482 3641
rect 517426 3567 517482 3576
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 518360 480 518388 3538
rect 519004 3466 519032 3703
rect 518992 3460 519044 3466
rect 518992 3402 519044 3408
rect 519556 480 519584 4150
rect 520752 480 520780 5782
rect 523040 4276 523092 4282
rect 523040 4218 523092 4224
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 521856 480 521884 3470
rect 523052 480 523080 4218
rect 524248 480 524276 5850
rect 526628 4480 526680 4486
rect 526628 4422 526680 4428
rect 525432 2644 525484 2650
rect 525432 2586 525484 2592
rect 525444 480 525472 2586
rect 526640 480 526668 4422
rect 527836 480 527864 6054
rect 530124 4548 530176 4554
rect 530124 4490 530176 4496
rect 529020 2848 529072 2854
rect 529020 2790 529072 2796
rect 529032 480 529060 2790
rect 530136 480 530164 4490
rect 531332 480 531360 6802
rect 534908 6792 534960 6798
rect 534908 6734 534960 6740
rect 533712 4616 533764 4622
rect 533712 4558 533764 4564
rect 532516 2916 532568 2922
rect 532516 2858 532568 2864
rect 532528 480 532556 2858
rect 533724 480 533752 4558
rect 534920 480 534948 6734
rect 538404 6724 538456 6730
rect 538404 6666 538456 6672
rect 537208 4684 537260 4690
rect 537208 4626 537260 4632
rect 536104 2984 536156 2990
rect 536104 2926 536156 2932
rect 536116 480 536144 2926
rect 537220 480 537248 4626
rect 538416 480 538444 6666
rect 541992 6656 542044 6662
rect 541992 6598 542044 6604
rect 540796 4752 540848 4758
rect 540796 4694 540848 4700
rect 539600 3052 539652 3058
rect 539600 2994 539652 3000
rect 539612 480 539640 2994
rect 540808 480 540836 4694
rect 542004 480 542032 6598
rect 545488 6452 545540 6458
rect 545488 6394 545540 6400
rect 544384 5364 544436 5370
rect 544384 5306 544436 5312
rect 543188 3120 543240 3126
rect 543188 3062 543240 3068
rect 543200 480 543228 3062
rect 544396 480 544424 5306
rect 545500 480 545528 6394
rect 549076 6384 549128 6390
rect 549076 6326 549128 6332
rect 547880 5296 547932 5302
rect 547880 5238 547932 5244
rect 546684 3188 546736 3194
rect 546684 3130 546736 3136
rect 546696 480 546724 3130
rect 547892 480 547920 5238
rect 549088 480 549116 6326
rect 552664 6316 552716 6322
rect 552664 6258 552716 6264
rect 551468 5228 551520 5234
rect 551468 5170 551520 5176
rect 550272 3392 550324 3398
rect 550272 3334 550324 3340
rect 550284 480 550312 3334
rect 551480 480 551508 5170
rect 552676 480 552704 6258
rect 556160 6248 556212 6254
rect 556160 6190 556212 6196
rect 554964 5160 555016 5166
rect 554964 5102 555016 5108
rect 553768 4140 553820 4146
rect 553768 4082 553820 4088
rect 553780 480 553808 4082
rect 554976 480 555004 5102
rect 556172 480 556200 6190
rect 559748 6180 559800 6186
rect 559748 6122 559800 6128
rect 558552 5092 558604 5098
rect 558552 5034 558604 5040
rect 557356 4072 557408 4078
rect 557356 4014 557408 4020
rect 557368 480 557396 4014
rect 558564 480 558592 5034
rect 559760 480 559788 6122
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 560864 480 560892 3946
rect 562060 480 562088 4966
rect 563256 480 563284 6938
rect 565636 4820 565688 4826
rect 565636 4762 565688 4768
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 564452 480 564480 3878
rect 565648 480 565676 4762
rect 566844 480 566872 7142
rect 568028 3732 568080 3738
rect 568028 3674 568080 3680
rect 568040 480 568068 3674
rect 569144 480 569172 16546
rect 570328 7268 570380 7274
rect 570328 7210 570380 7216
rect 570340 480 570368 7210
rect 571524 3664 571576 3670
rect 571524 3606 571576 3612
rect 571536 480 571564 3606
rect 572732 480 572760 77930
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 575480 35216 575532 35222
rect 575480 35158 575532 35164
rect 575492 16574 575520 35158
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20596 580224 20602
rect 580172 20538 580224 20544
rect 580184 19825 580212 20538
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 575492 16546 576348 16574
rect 573916 7336 573968 7342
rect 573916 7278 573968 7284
rect 573928 480 573956 7278
rect 575112 3596 575164 3602
rect 575112 3538 575164 3544
rect 575124 480 575152 3538
rect 576320 480 576348 16546
rect 577412 7472 577464 7478
rect 577412 7414 577464 7420
rect 577424 480 577452 7414
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580184 5846 580212 6559
rect 580172 5840 580224 5846
rect 580172 5782 580224 5788
rect 582194 3632 582250 3641
rect 582194 3567 582250 3576
rect 579804 3528 579856 3534
rect 578606 3496 578662 3505
rect 579804 3470 579856 3476
rect 578606 3431 578662 3440
rect 578620 480 578648 3431
rect 579816 480 579844 3470
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 3567
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 684256 3570 684312
rect 3422 671200 3478 671256
rect 580170 697176 580226 697232
rect 66994 679088 67050 679144
rect 580170 683848 580226 683904
rect 520922 678816 520978 678872
rect 67178 668888 67234 668944
rect 3514 658144 3570 658200
rect 67362 657736 67418 657792
rect 580170 670656 580226 670712
rect 521014 668480 521070 668536
rect 580170 657328 580226 657384
rect 520922 657192 520978 657248
rect 67362 646584 67418 646640
rect 521014 645768 521070 645824
rect 3422 645088 3478 645144
rect 580170 644000 580226 644056
rect 67362 635432 67418 635488
rect 520922 634480 520978 634536
rect 3422 632032 3478 632088
rect 580170 630808 580226 630864
rect 67362 624144 67418 624200
rect 520922 622920 520978 622976
rect 3422 619112 3478 619168
rect 580170 617480 580226 617536
rect 66902 612992 66958 613048
rect 520278 611632 520334 611688
rect 4066 606056 4122 606112
rect 580170 604152 580226 604208
rect 66442 601840 66498 601896
rect 521106 600208 521162 600264
rect 3422 593000 3478 593056
rect 579802 590960 579858 591016
rect 66994 590688 67050 590744
rect 521566 588784 521622 588840
rect 3422 579944 3478 580000
rect 67178 579572 67180 579592
rect 67180 579572 67232 579592
rect 67232 579572 67234 579592
rect 67178 579536 67234 579572
rect 580170 577632 580226 577688
rect 521566 577516 521622 577552
rect 521566 577496 521568 577516
rect 521568 577496 521620 577516
rect 521620 577496 521622 577516
rect 67362 568248 67418 568304
rect 4066 566888 4122 566944
rect 520738 566072 520794 566128
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 67362 557232 67418 557288
rect 521014 554648 521070 554704
rect 3422 553832 3478 553888
rect 579986 551112 580042 551168
rect 66626 545944 66682 546000
rect 520922 543224 520978 543280
rect 2962 540776 3018 540832
rect 580170 537784 580226 537840
rect 67362 534792 67418 534848
rect 520922 531936 520978 531992
rect 3422 527856 3478 527912
rect 579802 524456 579858 524512
rect 66442 523640 66498 523696
rect 520922 520512 520978 520568
rect 3422 514800 3478 514856
rect 67362 512352 67418 512408
rect 580170 511264 580226 511320
rect 521014 509088 521070 509144
rect 3422 501744 3478 501800
rect 67454 501336 67510 501392
rect 580170 497936 580226 497992
rect 520922 497800 520978 497856
rect 67454 490048 67510 490104
rect 3514 488688 3570 488744
rect 521014 486240 521070 486296
rect 67362 479032 67418 479088
rect 3422 475632 3478 475688
rect 520922 474952 520978 475008
rect 66994 467744 67050 467800
rect 3514 462576 3570 462632
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 521106 463528 521162 463584
rect 67362 456592 67418 456648
rect 3422 449520 3478 449576
rect 521014 452104 521070 452160
rect 66718 445440 66774 445496
rect 520922 440816 520978 440872
rect 3514 436600 3570 436656
rect 67178 434288 67234 434344
rect 3422 423544 3478 423600
rect 66810 423136 66866 423192
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 444760 580226 444816
rect 580170 431568 580226 431624
rect 521014 429392 521070 429448
rect 520922 418104 520978 418160
rect 67270 411848 67326 411904
rect 3606 410488 3662 410544
rect 67454 400832 67510 400888
rect 3514 397432 3570 397488
rect 3422 384376 3478 384432
rect 580170 418240 580226 418296
rect 521106 406680 521162 406736
rect 521014 395256 521070 395312
rect 67362 389544 67418 389600
rect 520922 383968 520978 384024
rect 67362 378392 67418 378448
rect 3606 371320 3662 371376
rect 67362 367240 67418 367296
rect 3514 358400 3570 358456
rect 3422 345344 3478 345400
rect 67362 356108 67418 356144
rect 67362 356088 67364 356108
rect 67364 356088 67416 356108
rect 67416 356088 67418 356108
rect 580170 404912 580226 404968
rect 580170 391720 580226 391776
rect 580170 378392 580226 378448
rect 521198 372408 521254 372464
rect 521106 361120 521162 361176
rect 521014 349832 521070 349888
rect 67362 344936 67418 344992
rect 520922 338272 520978 338328
rect 67178 333784 67234 333840
rect 3698 332288 3754 332344
rect 67362 322632 67418 322688
rect 3606 319232 3662 319288
rect 3514 306176 3570 306232
rect 3422 293120 3478 293176
rect 66718 311344 66774 311400
rect 67362 300192 67418 300248
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 338544 580226 338600
rect 521198 326984 521254 327040
rect 521106 315560 521162 315616
rect 521014 304136 521070 304192
rect 520922 292848 520978 292904
rect 66442 289040 66498 289096
rect 3698 280064 3754 280120
rect 67362 277888 67418 277944
rect 3606 267144 3662 267200
rect 3514 254088 3570 254144
rect 3422 241032 3478 241088
rect 67362 266736 67418 266792
rect 67362 255584 67418 255640
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 285368 580226 285424
rect 521290 281424 521346 281480
rect 521198 270000 521254 270056
rect 521106 258712 521162 258768
rect 521014 247288 521070 247344
rect 67362 244432 67418 244488
rect 520922 235864 520978 235920
rect 67178 233300 67234 233336
rect 67178 233280 67180 233300
rect 67180 233280 67232 233300
rect 67232 233280 67234 233300
rect 3790 227976 3846 228032
rect 67362 221992 67418 222048
rect 3698 214920 3754 214976
rect 3606 201864 3662 201920
rect 3514 188808 3570 188864
rect 3422 175888 3478 175944
rect 67362 210840 67418 210896
rect 67362 199688 67418 199744
rect 67454 188536 67510 188592
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 521382 224440 521438 224496
rect 521290 213152 521346 213208
rect 521198 201728 521254 201784
rect 521106 190304 521162 190360
rect 521014 179016 521070 179072
rect 67362 177384 67418 177440
rect 520922 167592 520978 167648
rect 67362 166232 67418 166288
rect 3882 162832 3938 162888
rect 67270 155080 67326 155136
rect 3790 149776 3846 149832
rect 3698 136720 3754 136776
rect 3606 123664 3662 123720
rect 3514 110608 3570 110664
rect 3422 97552 3478 97608
rect 67362 143792 67418 143848
rect 67178 132776 67234 132832
rect 67362 121508 67418 121544
rect 67362 121488 67364 121508
rect 67364 121488 67416 121508
rect 67416 121488 67418 121508
rect 67362 110336 67418 110392
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 521474 156168 521530 156224
rect 521382 144744 521438 144800
rect 521290 133456 521346 133512
rect 521198 122032 521254 122088
rect 521106 110608 521162 110664
rect 521014 99320 521070 99376
rect 67178 99184 67234 99240
rect 67454 89120 67510 89176
rect 520922 88848 520978 88904
rect 3974 84632 4030 84688
rect 3882 71576 3938 71632
rect 3790 58520 3846 58576
rect 3698 45464 3754 45520
rect 3606 32408 3662 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 11150 3440 11206 3496
rect 20626 3576 20682 3632
rect 25318 3712 25374 3768
rect 128358 2796 128360 2816
rect 128360 2796 128412 2816
rect 128412 2796 128414 2816
rect 128358 2760 128414 2796
rect 132222 2896 132278 2952
rect 132590 2760 132646 2816
rect 134062 2896 134118 2952
rect 160282 3440 160338 3496
rect 161570 3576 161626 3632
rect 162858 3712 162914 3768
rect 164330 3304 164386 3360
rect 205270 5244 205272 5264
rect 205272 5244 205324 5264
rect 205324 5244 205326 5264
rect 205270 5208 205326 5244
rect 205362 5072 205418 5128
rect 209686 5208 209742 5264
rect 209594 5072 209650 5128
rect 219438 5108 219440 5128
rect 219440 5108 219492 5128
rect 219492 5108 219494 5128
rect 219438 5072 219494 5108
rect 225142 5072 225198 5128
rect 248878 8880 248934 8936
rect 273258 9016 273314 9072
rect 273350 8916 273352 8936
rect 273352 8916 273404 8936
rect 273404 8916 273406 8936
rect 273350 8880 273406 8916
rect 277306 10376 277362 10432
rect 279514 10104 279570 10160
rect 282642 10920 282698 10976
rect 282826 10412 282828 10432
rect 282828 10412 282880 10432
rect 282880 10412 282882 10432
rect 282826 10376 282882 10412
rect 282918 9016 282974 9072
rect 292302 11092 292304 11112
rect 292304 11092 292356 11112
rect 292356 11092 292358 11112
rect 292302 11056 292358 11092
rect 292394 10104 292450 10160
rect 292394 9288 292450 9344
rect 292578 11192 292634 11248
rect 292578 10784 292634 10840
rect 292854 11192 292910 11248
rect 292946 11092 292948 11112
rect 292948 11092 293000 11112
rect 293000 11092 293002 11112
rect 292946 11056 293002 11092
rect 292946 9324 292948 9344
rect 292948 9324 293000 9344
rect 293000 9324 293002 9344
rect 292946 9288 293002 9324
rect 302330 10804 302386 10840
rect 302330 10784 302332 10804
rect 302332 10784 302384 10804
rect 302384 10784 302386 10804
rect 302330 10104 302386 10160
rect 302514 11076 302570 11112
rect 302514 11056 302516 11076
rect 302516 11056 302568 11076
rect 302568 11056 302570 11076
rect 311438 10376 311494 10432
rect 311714 10140 311716 10160
rect 311716 10140 311768 10160
rect 311768 10140 311770 10160
rect 311714 10104 311770 10140
rect 313462 10376 313518 10432
rect 316038 4936 316094 4992
rect 334162 4936 334218 4992
rect 348790 6604 348792 6624
rect 348792 6604 348844 6624
rect 348844 6604 348846 6624
rect 348790 6568 348846 6604
rect 354034 6568 354090 6624
rect 362314 3304 362370 3360
rect 369674 9152 369730 9208
rect 365810 3440 365866 3496
rect 369398 3576 369454 3632
rect 373906 9172 373962 9208
rect 373906 9152 373908 9172
rect 373908 9152 373960 9172
rect 373960 9152 373962 9172
rect 373722 9052 373724 9072
rect 373724 9052 373776 9072
rect 373776 9052 373778 9072
rect 373722 9016 373778 9052
rect 372894 3712 372950 3768
rect 383658 4936 383714 4992
rect 383658 4800 383714 4856
rect 393410 8916 393412 8936
rect 393412 8916 393464 8936
rect 393464 8916 393466 8936
rect 393410 8880 393466 8916
rect 393318 8744 393374 8800
rect 394514 6160 394570 6216
rect 398838 7112 398894 7168
rect 398654 6976 398710 7032
rect 398930 6996 398986 7032
rect 398930 6976 398932 6996
rect 398932 6976 398984 6996
rect 398984 6976 398986 6996
rect 403622 8744 403678 8800
rect 408314 7384 408370 7440
rect 408406 7148 408408 7168
rect 408408 7148 408460 7168
rect 408460 7148 408462 7168
rect 408406 7112 408462 7148
rect 412730 7420 412732 7440
rect 412732 7420 412784 7440
rect 412784 7420 412786 7440
rect 412730 7384 412786 7420
rect 412638 7248 412694 7304
rect 423770 7248 423826 7304
rect 441710 3848 441766 3904
rect 451278 3984 451334 4040
rect 451370 3884 451372 3904
rect 451372 3884 451424 3904
rect 451424 3884 451426 3904
rect 451370 3848 451426 3884
rect 454406 3848 454462 3904
rect 455510 3884 455512 3904
rect 455512 3884 455564 3904
rect 455564 3884 455566 3904
rect 455510 3848 455566 3884
rect 456798 3984 456854 4040
rect 458086 3848 458142 3904
rect 458178 3304 458234 3360
rect 459650 3576 459706 3632
rect 459742 3440 459798 3496
rect 460662 4120 460718 4176
rect 460570 4004 460626 4040
rect 460570 3984 460572 4004
rect 460572 3984 460624 4004
rect 460624 3984 460626 4004
rect 460846 3848 460902 3904
rect 461122 4020 461124 4040
rect 461124 4020 461176 4040
rect 461176 4020 461178 4040
rect 461122 3984 461178 4020
rect 460938 3712 460994 3768
rect 462318 4120 462374 4176
rect 460938 3032 460994 3088
rect 462318 3032 462374 3088
rect 463882 6196 463884 6216
rect 463884 6196 463936 6216
rect 463936 6196 463938 6216
rect 463882 6160 463938 6196
rect 470690 4800 470746 4856
rect 480350 4936 480406 4992
rect 480258 4820 480314 4856
rect 480258 4800 480260 4820
rect 480260 4800 480312 4820
rect 480312 4800 480314 4820
rect 489918 5072 489974 5128
rect 489826 4936 489882 4992
rect 499670 5516 499672 5536
rect 499672 5516 499724 5536
rect 499724 5516 499726 5536
rect 499670 5480 499726 5516
rect 499394 4936 499450 4992
rect 499762 4936 499818 4992
rect 499486 4820 499542 4856
rect 499486 4800 499488 4820
rect 499488 4800 499540 4820
rect 499540 4800 499542 4820
rect 506478 5480 506534 5536
rect 509238 4972 509240 4992
rect 509240 4972 509292 4992
rect 509292 4972 509294 4992
rect 509238 4936 509294 4972
rect 512458 4936 512514 4992
rect 511906 3848 511962 3904
rect 513286 3712 513342 3768
rect 514666 3440 514722 3496
rect 515862 3304 515918 3360
rect 516230 3732 516286 3768
rect 516230 3712 516232 3732
rect 516232 3712 516284 3732
rect 516284 3712 516286 3732
rect 518622 3848 518678 3904
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 518806 3712 518862 3768
rect 518990 3712 519046 3768
rect 517426 3576 517482 3632
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580170 6568 580226 6624
rect 582194 3576 582250 3632
rect 578606 3440 578662 3496
rect 580998 3304 581054 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 66989 679146 67055 679149
rect 66989 679144 69490 679146
rect 66989 679088 66994 679144
rect 67050 679140 69490 679144
rect 67050 679088 70012 679140
rect 66989 679086 70012 679088
rect 66989 679083 67055 679086
rect 69430 679080 70012 679086
rect 517868 678874 518450 678896
rect 520917 678874 520983 678877
rect 517868 678872 520983 678874
rect 517868 678836 520922 678872
rect 518390 678816 520922 678836
rect 520978 678816 520983 678872
rect 518390 678814 520983 678816
rect 520917 678811 520983 678814
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 67173 668946 67239 668949
rect 67173 668944 69490 668946
rect 67173 668888 67178 668944
rect 67234 668892 69490 668944
rect 67234 668888 70012 668892
rect 67173 668886 70012 668888
rect 67173 668883 67239 668886
rect 69430 668832 70012 668886
rect 521009 668538 521075 668541
rect 518390 668536 521075 668538
rect 518390 668526 521014 668536
rect 517868 668480 521014 668526
rect 521070 668480 521075 668536
rect 517868 668478 521075 668480
rect 517868 668466 518450 668478
rect 521009 668475 521075 668478
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 67357 657794 67423 657797
rect 67357 657792 69490 657794
rect 67357 657736 67362 657792
rect 67418 657790 69490 657792
rect 67418 657736 70012 657790
rect 67357 657734 70012 657736
rect 67357 657731 67423 657734
rect 69430 657730 70012 657734
rect 580165 657386 580231 657389
rect 583520 657386 584960 657476
rect 580165 657384 584960 657386
rect 580165 657328 580170 657384
rect 580226 657328 584960 657384
rect 580165 657326 584960 657328
rect 580165 657323 580231 657326
rect 520917 657250 520983 657253
rect 518390 657248 520983 657250
rect 518390 657192 520922 657248
rect 520978 657192 520983 657248
rect 583520 657236 584960 657326
rect 518390 657190 520983 657192
rect 518390 657180 518450 657190
rect 520917 657187 520983 657190
rect 517868 657120 518450 657180
rect 67357 646642 67423 646645
rect 67357 646640 69490 646642
rect 67357 646584 67362 646640
rect 67418 646584 69490 646640
rect 67357 646582 69490 646584
rect 67357 646579 67423 646582
rect 69430 646566 69490 646582
rect 69430 646506 70012 646566
rect 517868 645826 518450 645834
rect 521009 645826 521075 645829
rect 517868 645824 521075 645826
rect 517868 645774 521014 645824
rect 518390 645768 521014 645774
rect 521070 645768 521075 645824
rect 518390 645766 521075 645768
rect 521009 645763 521075 645766
rect -960 645146 480 645236
rect 3417 645146 3483 645149
rect -960 645144 3483 645146
rect -960 645088 3422 645144
rect 3478 645088 3483 645144
rect -960 645086 3483 645088
rect -960 644996 480 645086
rect 3417 645083 3483 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 67357 635490 67423 635493
rect 67357 635488 69490 635490
rect 67357 635432 67362 635488
rect 67418 635464 69490 635488
rect 67418 635432 70012 635464
rect 67357 635430 70012 635432
rect 67357 635427 67423 635430
rect 69430 635404 70012 635430
rect 520917 634538 520983 634541
rect 518390 634536 520983 634538
rect 518390 634488 520922 634536
rect 517868 634480 520922 634488
rect 520978 634480 520983 634536
rect 517868 634478 520983 634480
rect 517868 634428 518450 634478
rect 520917 634475 520983 634478
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 67357 624202 67423 624205
rect 69430 624202 70012 624240
rect 67357 624200 70012 624202
rect 67357 624144 67362 624200
rect 67418 624180 70012 624200
rect 67418 624144 69490 624180
rect 67357 624142 69490 624144
rect 67357 624139 67423 624142
rect 517868 622978 518450 623020
rect 520917 622978 520983 622981
rect 517868 622976 520983 622978
rect 517868 622960 520922 622976
rect 518390 622920 520922 622960
rect 520978 622920 520983 622976
rect 518390 622918 520983 622920
rect 520917 622915 520983 622918
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 66897 613050 66963 613053
rect 66897 613048 69490 613050
rect 66897 612992 66902 613048
rect 66958 613016 69490 613048
rect 66958 612992 70012 613016
rect 66897 612990 70012 612992
rect 66897 612987 66963 612990
rect 69430 612956 70012 612990
rect 520273 611690 520339 611693
rect 518390 611688 520339 611690
rect 518390 611674 520278 611688
rect 517868 611632 520278 611674
rect 520334 611632 520339 611688
rect 517868 611630 520339 611632
rect 517868 611614 518450 611630
rect 520273 611627 520339 611630
rect -960 606114 480 606204
rect 4061 606114 4127 606117
rect -960 606112 4127 606114
rect -960 606056 4066 606112
rect 4122 606056 4127 606112
rect -960 606054 4127 606056
rect -960 605964 480 606054
rect 4061 606051 4127 606054
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 66437 601898 66503 601901
rect 69430 601898 70012 601914
rect 66437 601896 70012 601898
rect 66437 601840 66442 601896
rect 66498 601854 70012 601896
rect 66498 601840 69490 601854
rect 66437 601838 69490 601840
rect 66437 601835 66503 601838
rect 517868 600268 518450 600328
rect 518390 600266 518450 600268
rect 521101 600266 521167 600269
rect 518390 600264 521167 600266
rect 518390 600208 521106 600264
rect 521162 600208 521167 600264
rect 518390 600206 521167 600208
rect 521101 600203 521167 600206
rect -960 593058 480 593148
rect 3417 593058 3483 593061
rect -960 593056 3483 593058
rect -960 593000 3422 593056
rect 3478 593000 3483 593056
rect -960 592998 3483 593000
rect -960 592908 480 592998
rect 3417 592995 3483 592998
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 66989 590746 67055 590749
rect 66989 590744 69490 590746
rect 66989 590688 66994 590744
rect 67050 590690 69490 590744
rect 67050 590688 70012 590690
rect 66989 590686 70012 590688
rect 66989 590683 67055 590686
rect 69430 590630 70012 590686
rect 517868 588842 518450 588860
rect 521561 588842 521627 588845
rect 517868 588840 521627 588842
rect 517868 588800 521566 588840
rect 518390 588784 521566 588800
rect 521622 588784 521627 588840
rect 518390 588782 521627 588784
rect 521561 588779 521627 588782
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 67173 579594 67239 579597
rect 67173 579592 69490 579594
rect 67173 579536 67178 579592
rect 67234 579588 69490 579592
rect 67234 579536 70012 579588
rect 67173 579534 70012 579536
rect 67173 579531 67239 579534
rect 69430 579528 70012 579534
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 521561 577554 521627 577557
rect 518390 577552 521627 577554
rect 518390 577514 521566 577552
rect 517868 577496 521566 577514
rect 521622 577496 521627 577552
rect 583520 577540 584960 577630
rect 517868 577494 521627 577496
rect 517868 577454 518450 577494
rect 521561 577491 521627 577494
rect 67357 568306 67423 568309
rect 69430 568306 70012 568364
rect 67357 568304 70012 568306
rect 67357 568248 67362 568304
rect 67418 568248 69490 568304
rect 67357 568246 69490 568248
rect 67357 568243 67423 568246
rect -960 566946 480 567036
rect 4061 566946 4127 566949
rect -960 566944 4127 566946
rect -960 566888 4066 566944
rect 4122 566888 4127 566944
rect -960 566886 4127 566888
rect -960 566796 480 566886
rect 4061 566883 4127 566886
rect 517868 566130 518450 566168
rect 520733 566130 520799 566133
rect 517868 566128 520799 566130
rect 517868 566108 520738 566128
rect 518390 566072 520738 566108
rect 520794 566072 520799 566128
rect 518390 566070 520799 566072
rect 520733 566067 520799 566070
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 67357 557290 67423 557293
rect 67357 557288 69490 557290
rect 67357 557232 67362 557288
rect 67418 557262 69490 557288
rect 67418 557232 70012 557262
rect 67357 557230 70012 557232
rect 67357 557227 67423 557230
rect 69430 557202 70012 557230
rect 521009 554706 521075 554709
rect 518390 554704 521075 554706
rect 518390 554700 521014 554704
rect 517868 554648 521014 554700
rect 521070 554648 521075 554704
rect 517868 554646 521075 554648
rect 517868 554640 518450 554646
rect 521009 554643 521075 554646
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 579981 551170 580047 551173
rect 583520 551170 584960 551260
rect 579981 551168 584960 551170
rect 579981 551112 579986 551168
rect 580042 551112 584960 551168
rect 579981 551110 584960 551112
rect 579981 551107 580047 551110
rect 583520 551020 584960 551110
rect 66621 546002 66687 546005
rect 69430 546002 70012 546038
rect 66621 546000 70012 546002
rect 66621 545944 66626 546000
rect 66682 545978 70012 546000
rect 66682 545944 69490 545978
rect 66621 545942 69490 545944
rect 66621 545939 66687 545942
rect 517868 543294 518450 543354
rect 518390 543282 518450 543294
rect 520917 543282 520983 543285
rect 518390 543280 520983 543282
rect 518390 543224 520922 543280
rect 520978 543224 520983 543280
rect 518390 543222 520983 543224
rect 520917 543219 520983 543222
rect -960 540834 480 540924
rect 2957 540834 3023 540837
rect -960 540832 3023 540834
rect -960 540776 2962 540832
rect 3018 540776 3023 540832
rect -960 540774 3023 540776
rect -960 540684 480 540774
rect 2957 540771 3023 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 69430 534876 70012 534936
rect 67357 534850 67423 534853
rect 69430 534850 69490 534876
rect 67357 534848 69490 534850
rect 67357 534792 67362 534848
rect 67418 534792 69490 534848
rect 67357 534790 69490 534792
rect 67357 534787 67423 534790
rect 517868 531994 518450 532008
rect 520917 531994 520983 531997
rect 517868 531992 520983 531994
rect 517868 531948 520922 531992
rect 518390 531936 520922 531948
rect 520978 531936 520983 531992
rect 518390 531934 520983 531936
rect 520917 531931 520983 531934
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect 66437 523698 66503 523701
rect 69430 523698 70012 523712
rect 66437 523696 70012 523698
rect 66437 523640 66442 523696
rect 66498 523652 70012 523696
rect 66498 523640 69490 523652
rect 66437 523638 69490 523640
rect 66437 523635 66503 523638
rect 520917 520570 520983 520573
rect 518390 520568 520983 520570
rect 518390 520540 520922 520568
rect 517868 520512 520922 520540
rect 520978 520512 520983 520568
rect 517868 520510 520983 520512
rect 517868 520480 518450 520510
rect 520917 520507 520983 520510
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 69430 512428 70012 512488
rect 67357 512410 67423 512413
rect 69430 512410 69490 512428
rect 67357 512408 69490 512410
rect 67357 512352 67362 512408
rect 67418 512352 69490 512408
rect 67357 512350 69490 512352
rect 67357 512347 67423 512350
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 517868 509146 518450 509194
rect 521009 509146 521075 509149
rect 517868 509144 521075 509146
rect 517868 509134 521014 509144
rect 518390 509088 521014 509134
rect 521070 509088 521075 509144
rect 518390 509086 521075 509088
rect 521009 509083 521075 509086
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 67449 501394 67515 501397
rect 67449 501392 69490 501394
rect 67449 501336 67454 501392
rect 67510 501386 69490 501392
rect 67510 501336 70012 501386
rect 67449 501334 70012 501336
rect 67449 501331 67515 501334
rect 69430 501326 70012 501334
rect 580165 497994 580231 497997
rect 583520 497994 584960 498084
rect 580165 497992 584960 497994
rect 580165 497936 580170 497992
rect 580226 497936 584960 497992
rect 580165 497934 584960 497936
rect 580165 497931 580231 497934
rect 520917 497858 520983 497861
rect 518390 497856 520983 497858
rect 518390 497848 520922 497856
rect 517868 497800 520922 497848
rect 520978 497800 520983 497856
rect 583520 497844 584960 497934
rect 517868 497798 520983 497800
rect 517868 497788 518450 497798
rect 520917 497795 520983 497798
rect 67449 490106 67515 490109
rect 69430 490106 70012 490162
rect 67449 490104 70012 490106
rect 67449 490048 67454 490104
rect 67510 490102 70012 490104
rect 67510 490048 69490 490102
rect 67449 490046 69490 490048
rect 67449 490043 67515 490046
rect -960 488746 480 488836
rect 3509 488746 3575 488749
rect -960 488744 3575 488746
rect -960 488688 3514 488744
rect 3570 488688 3575 488744
rect -960 488686 3575 488688
rect -960 488596 480 488686
rect 3509 488683 3575 488686
rect 517868 486320 518450 486380
rect 518390 486298 518450 486320
rect 521009 486298 521075 486301
rect 518390 486296 521075 486298
rect 518390 486240 521014 486296
rect 521070 486240 521075 486296
rect 518390 486238 521075 486240
rect 521009 486235 521075 486238
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 67357 479090 67423 479093
rect 67357 479088 69490 479090
rect 67357 479032 67362 479088
rect 67418 479060 69490 479088
rect 67418 479032 70012 479060
rect 67357 479030 70012 479032
rect 67357 479027 67423 479030
rect 69430 479000 70012 479030
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 517868 475010 518450 475034
rect 520917 475010 520983 475013
rect 517868 475008 520983 475010
rect 517868 474974 520922 475008
rect 518390 474952 520922 474974
rect 520978 474952 520983 475008
rect 518390 474950 520983 474952
rect 520917 474947 520983 474950
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 66989 467802 67055 467805
rect 69430 467802 70012 467836
rect 66989 467800 70012 467802
rect 66989 467744 66994 467800
rect 67050 467776 70012 467800
rect 67050 467744 69490 467776
rect 66989 467742 69490 467744
rect 66989 467739 67055 467742
rect 517868 463628 518450 463688
rect 518390 463586 518450 463628
rect 521101 463586 521167 463589
rect 518390 463584 521167 463586
rect 518390 463528 521106 463584
rect 521162 463528 521167 463584
rect 518390 463526 521167 463528
rect 521101 463523 521167 463526
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 69430 456674 70012 456734
rect 67357 456650 67423 456653
rect 69430 456650 69490 456674
rect 67357 456648 69490 456650
rect 67357 456592 67362 456648
rect 67418 456592 69490 456648
rect 67357 456590 69490 456592
rect 67357 456587 67423 456590
rect 517868 452162 518450 452220
rect 521009 452162 521075 452165
rect 517868 452160 521075 452162
rect 518390 452104 521014 452160
rect 521070 452104 521075 452160
rect 518390 452102 521075 452104
rect 521009 452099 521075 452102
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 66713 445498 66779 445501
rect 69430 445498 70012 445510
rect 66713 445496 70012 445498
rect 66713 445440 66718 445496
rect 66774 445450 70012 445496
rect 66774 445440 69490 445450
rect 66713 445438 69490 445440
rect 66713 445435 66779 445438
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 520917 440874 520983 440877
rect 517868 440872 520983 440874
rect 517868 440816 520922 440872
rect 520978 440816 520983 440872
rect 517868 440814 520983 440816
rect 520917 440811 520983 440814
rect -960 436658 480 436748
rect 3509 436658 3575 436661
rect -960 436656 3575 436658
rect -960 436600 3514 436656
rect 3570 436600 3575 436656
rect -960 436598 3575 436600
rect -960 436508 480 436598
rect 3509 436595 3575 436598
rect 67173 434346 67239 434349
rect 69430 434348 70012 434408
rect 69430 434346 69490 434348
rect 67173 434344 69490 434346
rect 67173 434288 67178 434344
rect 67234 434288 69490 434344
rect 67173 434286 69490 434288
rect 67173 434283 67239 434286
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 517868 429468 518450 429528
rect 518390 429450 518450 429468
rect 521009 429450 521075 429453
rect 518390 429448 521075 429450
rect 518390 429392 521014 429448
rect 521070 429392 521075 429448
rect 518390 429390 521075 429392
rect 521009 429387 521075 429390
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 66805 423194 66871 423197
rect 66805 423192 69490 423194
rect 66805 423136 66810 423192
rect 66866 423184 69490 423192
rect 66866 423136 70012 423184
rect 66805 423134 70012 423136
rect 66805 423131 66871 423134
rect 69430 423124 70012 423134
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 517868 418162 518082 418182
rect 520917 418162 520983 418165
rect 517868 418160 520983 418162
rect 517868 418122 520922 418160
rect 518022 418104 520922 418122
rect 520978 418104 520983 418160
rect 583520 418148 584960 418238
rect 518022 418102 520983 418104
rect 520917 418099 520983 418102
rect 67265 411906 67331 411909
rect 69430 411906 70012 411960
rect 67265 411904 70012 411906
rect 67265 411848 67270 411904
rect 67326 411900 70012 411904
rect 67326 411848 69490 411900
rect 67265 411846 69490 411848
rect 67265 411843 67331 411846
rect -960 410546 480 410636
rect 3601 410546 3667 410549
rect -960 410544 3667 410546
rect -960 410488 3606 410544
rect 3662 410488 3667 410544
rect -960 410486 3667 410488
rect -960 410396 480 410486
rect 3601 410483 3667 410486
rect 521101 406738 521167 406741
rect 518390 406736 521167 406738
rect 518390 406714 521106 406736
rect 517868 406680 521106 406714
rect 521162 406680 521167 406736
rect 517868 406678 521167 406680
rect 517868 406654 518450 406678
rect 521101 406675 521167 406678
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 67449 400890 67515 400893
rect 67449 400888 69490 400890
rect 67449 400832 67454 400888
rect 67510 400858 69490 400888
rect 67510 400832 70012 400858
rect 67449 400830 70012 400832
rect 67449 400827 67515 400830
rect 69430 400798 70012 400830
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 517868 395314 518450 395368
rect 521009 395314 521075 395317
rect 517868 395312 521075 395314
rect 517868 395308 521014 395312
rect 518390 395256 521014 395308
rect 521070 395256 521075 395312
rect 518390 395254 521075 395256
rect 521009 395251 521075 395254
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect 67357 389602 67423 389605
rect 69430 389602 70012 389634
rect 67357 389600 70012 389602
rect 67357 389544 67362 389600
rect 67418 389574 70012 389600
rect 67418 389544 69490 389574
rect 67357 389542 69490 389544
rect 67357 389539 67423 389542
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 520917 384026 520983 384029
rect 518390 384024 520983 384026
rect 518390 384022 520922 384024
rect 517868 383968 520922 384022
rect 520978 383968 520983 384024
rect 517868 383966 520983 383968
rect 517868 383962 518450 383966
rect 520917 383963 520983 383966
rect 69430 378472 70012 378532
rect 67357 378450 67423 378453
rect 69430 378450 69490 378472
rect 67357 378448 69490 378450
rect 67357 378392 67362 378448
rect 67418 378392 69490 378448
rect 67357 378390 69490 378392
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 67357 378387 67423 378390
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 517868 372494 518450 372554
rect 518390 372466 518450 372494
rect 521193 372466 521259 372469
rect 518390 372464 521259 372466
rect 518390 372408 521198 372464
rect 521254 372408 521259 372464
rect 518390 372406 521259 372408
rect 521193 372403 521259 372406
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 67357 367298 67423 367301
rect 69430 367298 70012 367308
rect 67357 367296 70012 367298
rect 67357 367240 67362 367296
rect 67418 367248 70012 367296
rect 67418 367240 69490 367248
rect 67357 367238 69490 367240
rect 67357 367235 67423 367238
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 517868 361178 518450 361208
rect 521101 361178 521167 361181
rect 517868 361176 521167 361178
rect 517868 361148 521106 361176
rect 518390 361120 521106 361148
rect 521162 361120 521167 361176
rect 518390 361118 521167 361120
rect 521101 361115 521167 361118
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 67357 356146 67423 356149
rect 69430 356146 70012 356206
rect 67357 356144 69490 356146
rect 67357 356088 67362 356144
rect 67418 356088 69490 356144
rect 67357 356086 69490 356088
rect 67357 356083 67423 356086
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 521009 349890 521075 349893
rect 518390 349888 521075 349890
rect 518390 349862 521014 349888
rect 517868 349832 521014 349862
rect 521070 349832 521075 349888
rect 517868 349830 521075 349832
rect 517868 349802 518450 349830
rect 521009 349827 521075 349830
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 67357 344994 67423 344997
rect 67357 344992 69490 344994
rect 67357 344936 67362 344992
rect 67418 344982 69490 344992
rect 67418 344936 70012 344982
rect 67357 344934 70012 344936
rect 67357 344931 67423 344934
rect 69430 344922 70012 344934
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 580165 338600 584960 338602
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect 517868 338334 518450 338394
rect 518390 338330 518450 338334
rect 520917 338330 520983 338333
rect 518390 338328 520983 338330
rect 518390 338272 520922 338328
rect 520978 338272 520983 338328
rect 518390 338270 520983 338272
rect 520917 338267 520983 338270
rect 67173 333842 67239 333845
rect 69430 333842 70012 333880
rect 67173 333840 70012 333842
rect 67173 333784 67178 333840
rect 67234 333820 70012 333840
rect 67234 333784 69490 333820
rect 67173 333782 69490 333784
rect 67173 333779 67239 333782
rect -960 332346 480 332436
rect 3693 332346 3759 332349
rect -960 332344 3759 332346
rect -960 332288 3698 332344
rect 3754 332288 3759 332344
rect -960 332286 3759 332288
rect -960 332196 480 332286
rect 3693 332283 3759 332286
rect 517868 327042 518450 327048
rect 521193 327042 521259 327045
rect 517868 327040 521259 327042
rect 517868 326988 521198 327040
rect 518390 326984 521198 326988
rect 521254 326984 521259 327040
rect 518390 326982 521259 326984
rect 521193 326979 521259 326982
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 67357 322690 67423 322693
rect 67357 322688 69490 322690
rect 67357 322632 67362 322688
rect 67418 322656 69490 322688
rect 67418 322632 70012 322656
rect 67357 322630 70012 322632
rect 67357 322627 67423 322630
rect 69430 322596 70012 322630
rect -960 319290 480 319380
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 517868 315642 518450 315702
rect 518390 315618 518450 315642
rect 521101 315618 521167 315621
rect 518390 315616 521167 315618
rect 518390 315560 521106 315616
rect 521162 315560 521167 315616
rect 518390 315558 521167 315560
rect 521101 315555 521167 315558
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 66713 311402 66779 311405
rect 69430 311402 70012 311432
rect 66713 311400 70012 311402
rect 66713 311344 66718 311400
rect 66774 311372 70012 311400
rect 66774 311344 69490 311372
rect 66713 311342 69490 311344
rect 66713 311339 66779 311342
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 517868 304194 518450 304234
rect 521009 304194 521075 304197
rect 517868 304192 521075 304194
rect 517868 304174 521014 304192
rect 518390 304136 521014 304174
rect 521070 304136 521075 304192
rect 518390 304134 521075 304136
rect 521009 304131 521075 304134
rect 69430 300270 70012 300330
rect 67357 300250 67423 300253
rect 69430 300250 69490 300270
rect 67357 300248 69490 300250
rect 67357 300192 67362 300248
rect 67418 300192 69490 300248
rect 67357 300190 69490 300192
rect 67357 300187 67423 300190
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 520917 292906 520983 292909
rect 518390 292904 520983 292906
rect 518390 292888 520922 292904
rect 517868 292848 520922 292888
rect 520978 292848 520983 292904
rect 517868 292846 520983 292848
rect 517868 292828 518450 292846
rect 520917 292843 520983 292846
rect 66437 289098 66503 289101
rect 69430 289098 70012 289106
rect 66437 289096 70012 289098
rect 66437 289040 66442 289096
rect 66498 289046 70012 289096
rect 66498 289040 69490 289046
rect 66437 289038 69490 289040
rect 66437 289035 66503 289038
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 517868 281482 518450 281542
rect 521285 281482 521351 281485
rect 518390 281480 521351 281482
rect 518390 281424 521290 281480
rect 521346 281424 521351 281480
rect 518390 281422 521351 281424
rect 521285 281419 521351 281422
rect -960 280122 480 280212
rect 3693 280122 3759 280125
rect -960 280120 3759 280122
rect -960 280064 3698 280120
rect 3754 280064 3759 280120
rect -960 280062 3759 280064
rect -960 279972 480 280062
rect 3693 280059 3759 280062
rect 67357 277946 67423 277949
rect 69430 277946 70012 278004
rect 67357 277944 70012 277946
rect 67357 277888 67362 277944
rect 67418 277888 69490 277944
rect 67357 277886 69490 277888
rect 67357 277883 67423 277886
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 517868 270058 518450 270074
rect 521193 270058 521259 270061
rect 517868 270056 521259 270058
rect 517868 270014 521198 270056
rect 518390 270000 521198 270014
rect 521254 270000 521259 270056
rect 518390 269998 521259 270000
rect 521193 269995 521259 269998
rect -960 267202 480 267292
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 67357 266794 67423 266797
rect 67357 266792 69490 266794
rect 67357 266736 67362 266792
rect 67418 266780 69490 266792
rect 67418 266736 70012 266780
rect 67357 266734 70012 266736
rect 67357 266731 67423 266734
rect 69430 266720 70012 266734
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 521101 258770 521167 258773
rect 518390 258768 521167 258770
rect 518390 258728 521106 258768
rect 517868 258712 521106 258728
rect 521162 258712 521167 258768
rect 583520 258756 584960 258846
rect 517868 258710 521167 258712
rect 517868 258668 518450 258710
rect 521101 258707 521167 258710
rect 67357 255642 67423 255645
rect 69430 255642 70012 255678
rect 67357 255640 70012 255642
rect 67357 255584 67362 255640
rect 67418 255618 70012 255640
rect 67418 255584 69490 255618
rect 67357 255582 69490 255584
rect 67357 255579 67423 255582
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 517868 247346 518450 247382
rect 521009 247346 521075 247349
rect 517868 247344 521075 247346
rect 517868 247322 521014 247344
rect 518390 247288 521014 247322
rect 521070 247288 521075 247344
rect 518390 247286 521075 247288
rect 521009 247283 521075 247286
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 67357 244490 67423 244493
rect 67357 244488 69490 244490
rect 67357 244432 67362 244488
rect 67418 244454 69490 244488
rect 67418 244432 70012 244454
rect 67357 244430 70012 244432
rect 67357 244427 67423 244430
rect 69430 244394 70012 244430
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 520917 235922 520983 235925
rect 518390 235920 520983 235922
rect 518390 235914 520922 235920
rect 517868 235864 520922 235914
rect 520978 235864 520983 235920
rect 517868 235862 520983 235864
rect 517868 235854 518450 235862
rect 520917 235859 520983 235862
rect 67173 233338 67239 233341
rect 69430 233338 70012 233352
rect 67173 233336 70012 233338
rect 67173 233280 67178 233336
rect 67234 233292 70012 233336
rect 67234 233280 69490 233292
rect 67173 233278 69490 233280
rect 67173 233275 67239 233278
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3785 228034 3851 228037
rect -960 228032 3851 228034
rect -960 227976 3790 228032
rect 3846 227976 3851 228032
rect -960 227974 3851 227976
rect -960 227884 480 227974
rect 3785 227971 3851 227974
rect 517868 224508 518450 224568
rect 518390 224498 518450 224508
rect 521377 224498 521443 224501
rect 518390 224496 521443 224498
rect 518390 224440 521382 224496
rect 521438 224440 521443 224496
rect 518390 224438 521443 224440
rect 521377 224435 521443 224438
rect 69430 222068 70012 222128
rect 67357 222050 67423 222053
rect 69430 222050 69490 222068
rect 67357 222048 69490 222050
rect 67357 221992 67362 222048
rect 67418 221992 69490 222048
rect 67357 221990 69490 221992
rect 67357 221987 67423 221990
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3693 214978 3759 214981
rect -960 214976 3759 214978
rect -960 214920 3698 214976
rect 3754 214920 3759 214976
rect -960 214918 3759 214920
rect -960 214828 480 214918
rect 3693 214915 3759 214918
rect 517868 213210 518450 213222
rect 521285 213210 521351 213213
rect 517868 213208 521351 213210
rect 517868 213162 521290 213208
rect 518390 213152 521290 213162
rect 521346 213152 521351 213208
rect 518390 213150 521351 213152
rect 521285 213147 521351 213150
rect 67357 210898 67423 210901
rect 69430 210898 70012 210904
rect 67357 210896 70012 210898
rect 67357 210840 67362 210896
rect 67418 210844 70012 210896
rect 67418 210840 69490 210844
rect 67357 210838 69490 210840
rect 67357 210835 67423 210838
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 517868 201816 518450 201876
rect 518390 201786 518450 201816
rect 521193 201786 521259 201789
rect 518390 201784 521259 201786
rect 518390 201728 521198 201784
rect 521254 201728 521259 201784
rect 518390 201726 521259 201728
rect 521193 201723 521259 201726
rect 67357 199746 67423 199749
rect 69430 199746 70012 199802
rect 67357 199744 70012 199746
rect 67357 199688 67362 199744
rect 67418 199742 70012 199744
rect 67418 199688 69490 199742
rect 67357 199686 69490 199688
rect 67357 199683 67423 199686
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 517868 190362 518450 190408
rect 521101 190362 521167 190365
rect 517868 190360 521167 190362
rect 517868 190348 521106 190360
rect 518390 190304 521106 190348
rect 521162 190304 521167 190360
rect 518390 190302 521167 190304
rect 521101 190299 521167 190302
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 67449 188594 67515 188597
rect 67449 188592 69490 188594
rect 67449 188536 67454 188592
rect 67510 188578 69490 188592
rect 67510 188536 70012 188578
rect 67449 188534 70012 188536
rect 67449 188531 67515 188534
rect 69430 188518 70012 188534
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 521009 179074 521075 179077
rect 518390 179072 521075 179074
rect 518390 179062 521014 179072
rect 517868 179016 521014 179062
rect 521070 179016 521075 179072
rect 583520 179060 584960 179150
rect 517868 179014 521075 179016
rect 517868 179002 518450 179014
rect 521009 179011 521075 179014
rect 67357 177442 67423 177445
rect 69430 177442 70012 177476
rect 67357 177440 70012 177442
rect 67357 177384 67362 177440
rect 67418 177416 70012 177440
rect 67418 177384 69490 177416
rect 67357 177382 69490 177384
rect 67357 177379 67423 177382
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 517868 167656 518450 167716
rect 518390 167650 518450 167656
rect 520917 167650 520983 167653
rect 518390 167648 520983 167650
rect 518390 167592 520922 167648
rect 520978 167592 520983 167648
rect 518390 167590 520983 167592
rect 520917 167587 520983 167590
rect 67357 166290 67423 166293
rect 67357 166288 69490 166290
rect 67357 166232 67362 166288
rect 67418 166252 69490 166288
rect 67418 166232 70012 166252
rect 67357 166230 70012 166232
rect 67357 166227 67423 166230
rect 69430 166192 70012 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3877 162890 3943 162893
rect -960 162888 3943 162890
rect -960 162832 3882 162888
rect 3938 162832 3943 162888
rect -960 162830 3943 162832
rect -960 162740 480 162830
rect 3877 162827 3943 162830
rect 517868 156226 518450 156248
rect 521469 156226 521535 156229
rect 517868 156224 521535 156226
rect 517868 156188 521474 156224
rect 518390 156168 521474 156188
rect 521530 156168 521535 156224
rect 518390 156166 521535 156168
rect 521469 156163 521535 156166
rect 67265 155138 67331 155141
rect 69430 155138 70012 155150
rect 67265 155136 70012 155138
rect 67265 155080 67270 155136
rect 67326 155090 70012 155136
rect 67326 155080 69490 155090
rect 67265 155078 69490 155080
rect 67265 155075 67331 155078
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3785 149834 3851 149837
rect -960 149832 3851 149834
rect -960 149776 3790 149832
rect 3846 149776 3851 149832
rect -960 149774 3851 149776
rect -960 149684 480 149774
rect 3785 149771 3851 149774
rect 517868 144842 518450 144902
rect 518390 144802 518450 144842
rect 521377 144802 521443 144805
rect 518390 144800 521443 144802
rect 518390 144744 521382 144800
rect 521438 144744 521443 144800
rect 518390 144742 521443 144744
rect 521377 144739 521443 144742
rect 69430 143866 70012 143926
rect 67357 143850 67423 143853
rect 69430 143850 69490 143866
rect 67357 143848 69490 143850
rect 67357 143792 67362 143848
rect 67418 143792 69490 143848
rect 67357 143790 69490 143792
rect 67357 143787 67423 143790
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 517868 133514 518450 133556
rect 521285 133514 521351 133517
rect 517868 133512 521351 133514
rect 517868 133496 521290 133512
rect 518390 133456 521290 133496
rect 521346 133456 521351 133512
rect 518390 133454 521351 133456
rect 521285 133451 521351 133454
rect 67173 132834 67239 132837
rect 67173 132832 69490 132834
rect 67173 132776 67178 132832
rect 67234 132824 69490 132832
rect 67234 132776 70012 132824
rect 67173 132774 70012 132776
rect 67173 132771 67239 132774
rect 69430 132764 70012 132774
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3601 123722 3667 123725
rect -960 123720 3667 123722
rect -960 123664 3606 123720
rect 3662 123664 3667 123720
rect -960 123662 3667 123664
rect -960 123572 480 123662
rect 3601 123659 3667 123662
rect 521193 122090 521259 122093
rect 518390 122088 521259 122090
rect 517868 122032 521198 122088
rect 521254 122032 521259 122088
rect 517868 122030 521259 122032
rect 517868 122028 518450 122030
rect 521193 122027 521259 122030
rect 67357 121546 67423 121549
rect 69430 121546 70012 121600
rect 67357 121544 70012 121546
rect 67357 121488 67362 121544
rect 67418 121540 70012 121544
rect 67418 121488 69490 121540
rect 67357 121486 69490 121488
rect 67357 121483 67423 121486
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 517868 110682 518450 110742
rect 3509 110666 3575 110669
rect -960 110664 3575 110666
rect -960 110608 3514 110664
rect 3570 110608 3575 110664
rect -960 110606 3575 110608
rect 518390 110666 518450 110682
rect 521101 110666 521167 110669
rect 518390 110664 521167 110666
rect 518390 110608 521106 110664
rect 521162 110608 521167 110664
rect 518390 110606 521167 110608
rect -960 110516 480 110606
rect 3509 110603 3575 110606
rect 521101 110603 521167 110606
rect 67357 110394 67423 110397
rect 67357 110392 69490 110394
rect 67357 110336 67362 110392
rect 67418 110376 69490 110392
rect 67418 110336 70012 110376
rect 67357 110334 70012 110336
rect 67357 110331 67423 110334
rect 69430 110316 70012 110334
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 517868 99378 518082 99396
rect 521009 99378 521075 99381
rect 517868 99376 521075 99378
rect 517868 99336 521014 99376
rect 518022 99320 521014 99336
rect 521070 99320 521075 99376
rect 583520 99364 584960 99454
rect 518022 99318 521075 99320
rect 521009 99315 521075 99318
rect 67173 99242 67239 99245
rect 69430 99242 70012 99274
rect 67173 99240 70012 99242
rect 67173 99184 67178 99240
rect 67234 99214 70012 99240
rect 67234 99184 69490 99214
rect 67173 99182 69490 99184
rect 67173 99179 67239 99182
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 67449 89178 67515 89181
rect 67449 89176 69490 89178
rect 67449 89120 67454 89176
rect 67510 89148 69490 89176
rect 67510 89120 70012 89148
rect 67449 89118 70012 89120
rect 67449 89115 67515 89118
rect 69430 89088 70012 89118
rect 520917 88906 520983 88909
rect 518390 88904 520983 88906
rect 517868 88848 520922 88904
rect 520978 88848 520983 88904
rect 517868 88846 520983 88848
rect 517868 88844 518450 88846
rect 520917 88843 520983 88846
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3969 84690 4035 84693
rect -960 84688 4035 84690
rect -960 84632 3974 84688
rect 4030 84632 4035 84688
rect -960 84630 4035 84632
rect -960 84540 480 84630
rect 3969 84627 4035 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3877 71634 3943 71637
rect -960 71632 3943 71634
rect -960 71576 3882 71632
rect 3938 71576 3943 71632
rect -960 71574 3943 71576
rect -960 71484 480 71574
rect 3877 71571 3943 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3785 58578 3851 58581
rect -960 58576 3851 58578
rect -960 58520 3790 58576
rect 3846 58520 3851 58576
rect -960 58518 3851 58520
rect -960 58428 480 58518
rect 3785 58515 3851 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 292573 11250 292639 11253
rect 292849 11250 292915 11253
rect 292573 11248 292915 11250
rect 292573 11192 292578 11248
rect 292634 11192 292854 11248
rect 292910 11192 292915 11248
rect 292573 11190 292915 11192
rect 292573 11187 292639 11190
rect 292849 11187 292915 11190
rect 292297 11114 292363 11117
rect 292941 11114 293007 11117
rect 302509 11114 302575 11117
rect 292297 11112 293007 11114
rect 292297 11056 292302 11112
rect 292358 11056 292946 11112
rect 293002 11056 293007 11112
rect 292297 11054 293007 11056
rect 292297 11051 292363 11054
rect 292941 11051 293007 11054
rect 302190 11112 302575 11114
rect 302190 11056 302514 11112
rect 302570 11056 302575 11112
rect 302190 11054 302575 11056
rect 282637 10978 282703 10981
rect 302190 10978 302250 11054
rect 302509 11051 302575 11054
rect 282637 10976 302250 10978
rect 282637 10920 282642 10976
rect 282698 10920 302250 10976
rect 282637 10918 302250 10920
rect 282637 10915 282703 10918
rect 292573 10842 292639 10845
rect 302325 10842 302391 10845
rect 292573 10840 302391 10842
rect 292573 10784 292578 10840
rect 292634 10784 302330 10840
rect 302386 10784 302391 10840
rect 292573 10782 302391 10784
rect 292573 10779 292639 10782
rect 302325 10779 302391 10782
rect 277301 10434 277367 10437
rect 282821 10434 282887 10437
rect 277301 10432 282887 10434
rect 277301 10376 277306 10432
rect 277362 10376 282826 10432
rect 282882 10376 282887 10432
rect 277301 10374 282887 10376
rect 277301 10371 277367 10374
rect 282821 10371 282887 10374
rect 311433 10434 311499 10437
rect 313457 10434 313523 10437
rect 311433 10432 313523 10434
rect 311433 10376 311438 10432
rect 311494 10376 313462 10432
rect 313518 10376 313523 10432
rect 311433 10374 313523 10376
rect 311433 10371 311499 10374
rect 313457 10371 313523 10374
rect 279509 10162 279575 10165
rect 292389 10162 292455 10165
rect 279509 10160 292455 10162
rect 279509 10104 279514 10160
rect 279570 10104 292394 10160
rect 292450 10104 292455 10160
rect 279509 10102 292455 10104
rect 279509 10099 279575 10102
rect 292389 10099 292455 10102
rect 302325 10162 302391 10165
rect 311709 10162 311775 10165
rect 302325 10160 311775 10162
rect 302325 10104 302330 10160
rect 302386 10104 311714 10160
rect 311770 10104 311775 10160
rect 302325 10102 311775 10104
rect 302325 10099 302391 10102
rect 311709 10099 311775 10102
rect 292389 9346 292455 9349
rect 292941 9346 293007 9349
rect 292389 9344 293007 9346
rect 292389 9288 292394 9344
rect 292450 9288 292946 9344
rect 293002 9288 293007 9344
rect 292389 9286 293007 9288
rect 292389 9283 292455 9286
rect 292941 9283 293007 9286
rect 369669 9210 369735 9213
rect 373901 9210 373967 9213
rect 369669 9208 373967 9210
rect 369669 9152 369674 9208
rect 369730 9152 373906 9208
rect 373962 9152 373967 9208
rect 369669 9150 373967 9152
rect 369669 9147 369735 9150
rect 373901 9147 373967 9150
rect 273253 9074 273319 9077
rect 282913 9074 282979 9077
rect 273253 9072 282979 9074
rect 273253 9016 273258 9072
rect 273314 9016 282918 9072
rect 282974 9016 282979 9072
rect 273253 9014 282979 9016
rect 273253 9011 273319 9014
rect 282913 9011 282979 9014
rect 373717 9074 373783 9077
rect 373717 9072 383670 9074
rect 373717 9016 373722 9072
rect 373778 9016 383670 9072
rect 373717 9014 383670 9016
rect 373717 9011 373783 9014
rect 248873 8938 248939 8941
rect 273345 8938 273411 8941
rect 248873 8936 273411 8938
rect 248873 8880 248878 8936
rect 248934 8880 273350 8936
rect 273406 8880 273411 8936
rect 248873 8878 273411 8880
rect 383610 8938 383670 9014
rect 393405 8938 393471 8941
rect 383610 8936 393471 8938
rect 383610 8880 393410 8936
rect 393466 8880 393471 8936
rect 383610 8878 393471 8880
rect 248873 8875 248939 8878
rect 273345 8875 273411 8878
rect 393405 8875 393471 8878
rect 393313 8802 393379 8805
rect 403617 8802 403683 8805
rect 393313 8800 403683 8802
rect 393313 8744 393318 8800
rect 393374 8744 403622 8800
rect 403678 8744 403683 8800
rect 393313 8742 403683 8744
rect 393313 8739 393379 8742
rect 403617 8739 403683 8742
rect 408309 7442 408375 7445
rect 412725 7442 412791 7445
rect 408309 7440 412791 7442
rect 408309 7384 408314 7440
rect 408370 7384 412730 7440
rect 412786 7384 412791 7440
rect 408309 7382 412791 7384
rect 408309 7379 408375 7382
rect 412725 7379 412791 7382
rect 412633 7306 412699 7309
rect 423765 7306 423831 7309
rect 412633 7304 423831 7306
rect 412633 7248 412638 7304
rect 412694 7248 423770 7304
rect 423826 7248 423831 7304
rect 412633 7246 423831 7248
rect 412633 7243 412699 7246
rect 423765 7243 423831 7246
rect 398833 7170 398899 7173
rect 408401 7170 408467 7173
rect 398833 7168 408467 7170
rect 398833 7112 398838 7168
rect 398894 7112 408406 7168
rect 408462 7112 408467 7168
rect 398833 7110 408467 7112
rect 398833 7107 398899 7110
rect 408401 7107 408467 7110
rect 398649 7034 398715 7037
rect 398925 7034 398991 7037
rect 398649 7032 398991 7034
rect 398649 6976 398654 7032
rect 398710 6976 398930 7032
rect 398986 6976 398991 7032
rect 398649 6974 398991 6976
rect 398649 6971 398715 6974
rect 398925 6971 398991 6974
rect 348785 6626 348851 6629
rect 354029 6626 354095 6629
rect 348785 6624 354095 6626
rect -960 6490 480 6580
rect 348785 6568 348790 6624
rect 348846 6568 354034 6624
rect 354090 6568 354095 6624
rect 348785 6566 354095 6568
rect 348785 6563 348851 6566
rect 354029 6563 354095 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 394509 6218 394575 6221
rect 463877 6218 463943 6221
rect 394509 6216 463943 6218
rect 394509 6160 394514 6216
rect 394570 6160 463882 6216
rect 463938 6160 463943 6216
rect 394509 6158 463943 6160
rect 394509 6155 394575 6158
rect 463877 6155 463943 6158
rect 499665 5538 499731 5541
rect 506473 5538 506539 5541
rect 499665 5536 506539 5538
rect 499665 5480 499670 5536
rect 499726 5480 506478 5536
rect 506534 5480 506539 5536
rect 499665 5478 506539 5480
rect 499665 5475 499731 5478
rect 506473 5475 506539 5478
rect 205265 5266 205331 5269
rect 209681 5266 209747 5269
rect 205265 5264 209747 5266
rect 205265 5208 205270 5264
rect 205326 5208 209686 5264
rect 209742 5208 209747 5264
rect 205265 5206 209747 5208
rect 205265 5203 205331 5206
rect 209681 5203 209747 5206
rect 205357 5130 205423 5133
rect 209589 5130 209655 5133
rect 205357 5128 209655 5130
rect 205357 5072 205362 5128
rect 205418 5072 209594 5128
rect 209650 5072 209655 5128
rect 205357 5070 209655 5072
rect 205357 5067 205423 5070
rect 209589 5067 209655 5070
rect 219433 5130 219499 5133
rect 225137 5130 225203 5133
rect 489913 5130 489979 5133
rect 219433 5128 225203 5130
rect 219433 5072 219438 5128
rect 219494 5072 225142 5128
rect 225198 5072 225203 5128
rect 219433 5070 225203 5072
rect 219433 5067 219499 5070
rect 225137 5067 225203 5070
rect 489870 5128 489979 5130
rect 489870 5072 489918 5128
rect 489974 5072 489979 5128
rect 489870 5067 489979 5072
rect 489870 4997 489930 5067
rect 316033 4994 316099 4997
rect 334157 4994 334223 4997
rect 316033 4992 334223 4994
rect 316033 4936 316038 4992
rect 316094 4936 334162 4992
rect 334218 4936 334223 4992
rect 316033 4934 334223 4936
rect 316033 4931 316099 4934
rect 334157 4931 334223 4934
rect 383653 4994 383719 4997
rect 480345 4994 480411 4997
rect 383653 4992 480411 4994
rect 383653 4936 383658 4992
rect 383714 4936 480350 4992
rect 480406 4936 480411 4992
rect 383653 4934 480411 4936
rect 383653 4931 383719 4934
rect 480345 4931 480411 4934
rect 489821 4992 489930 4997
rect 489821 4936 489826 4992
rect 489882 4936 489930 4992
rect 489821 4934 489930 4936
rect 499389 4994 499455 4997
rect 499757 4994 499823 4997
rect 499389 4992 499823 4994
rect 499389 4936 499394 4992
rect 499450 4936 499762 4992
rect 499818 4936 499823 4992
rect 499389 4934 499823 4936
rect 489821 4931 489887 4934
rect 499389 4931 499455 4934
rect 499757 4931 499823 4934
rect 509233 4994 509299 4997
rect 512453 4994 512519 4997
rect 509233 4992 512519 4994
rect 509233 4936 509238 4992
rect 509294 4936 512458 4992
rect 512514 4936 512519 4992
rect 509233 4934 512519 4936
rect 509233 4931 509299 4934
rect 512453 4931 512519 4934
rect 383653 4858 383719 4861
rect 470685 4858 470751 4861
rect 383653 4856 470751 4858
rect 383653 4800 383658 4856
rect 383714 4800 470690 4856
rect 470746 4800 470751 4856
rect 383653 4798 470751 4800
rect 383653 4795 383719 4798
rect 470685 4795 470751 4798
rect 480253 4858 480319 4861
rect 499481 4858 499547 4861
rect 480253 4856 499547 4858
rect 480253 4800 480258 4856
rect 480314 4800 499486 4856
rect 499542 4800 499547 4856
rect 480253 4798 499547 4800
rect 480253 4795 480319 4798
rect 499481 4795 499547 4798
rect 460657 4178 460723 4181
rect 462313 4178 462379 4181
rect 460657 4176 462379 4178
rect 460657 4120 460662 4176
rect 460718 4120 462318 4176
rect 462374 4120 462379 4176
rect 460657 4118 462379 4120
rect 460657 4115 460723 4118
rect 462313 4115 462379 4118
rect 451273 4042 451339 4045
rect 456793 4042 456859 4045
rect 451273 4040 456859 4042
rect 451273 3984 451278 4040
rect 451334 3984 456798 4040
rect 456854 3984 456859 4040
rect 451273 3982 456859 3984
rect 451273 3979 451339 3982
rect 456793 3979 456859 3982
rect 460565 4042 460631 4045
rect 461117 4042 461183 4045
rect 460565 4040 461183 4042
rect 460565 3984 460570 4040
rect 460626 3984 461122 4040
rect 461178 3984 461183 4040
rect 460565 3982 461183 3984
rect 460565 3979 460631 3982
rect 461117 3979 461183 3982
rect 441705 3906 441771 3909
rect 451365 3906 451431 3909
rect 441705 3904 451431 3906
rect 441705 3848 441710 3904
rect 441766 3848 451370 3904
rect 451426 3848 451431 3904
rect 441705 3846 451431 3848
rect 441705 3843 441771 3846
rect 451365 3843 451431 3846
rect 454401 3906 454467 3909
rect 455505 3906 455571 3909
rect 454401 3904 455571 3906
rect 454401 3848 454406 3904
rect 454462 3848 455510 3904
rect 455566 3848 455571 3904
rect 454401 3846 455571 3848
rect 454401 3843 454467 3846
rect 455505 3843 455571 3846
rect 458081 3906 458147 3909
rect 460841 3906 460907 3909
rect 458081 3904 460907 3906
rect 458081 3848 458086 3904
rect 458142 3848 460846 3904
rect 460902 3848 460907 3904
rect 458081 3846 460907 3848
rect 458081 3843 458147 3846
rect 460841 3843 460907 3846
rect 511901 3906 511967 3909
rect 518617 3906 518683 3909
rect 511901 3904 518683 3906
rect 511901 3848 511906 3904
rect 511962 3848 518622 3904
rect 518678 3848 518683 3904
rect 511901 3846 518683 3848
rect 511901 3843 511967 3846
rect 518617 3843 518683 3846
rect 25313 3770 25379 3773
rect 162853 3770 162919 3773
rect 25313 3768 162919 3770
rect 25313 3712 25318 3768
rect 25374 3712 162858 3768
rect 162914 3712 162919 3768
rect 25313 3710 162919 3712
rect 25313 3707 25379 3710
rect 162853 3707 162919 3710
rect 372889 3770 372955 3773
rect 460933 3770 460999 3773
rect 372889 3768 460999 3770
rect 372889 3712 372894 3768
rect 372950 3712 460938 3768
rect 460994 3712 460999 3768
rect 372889 3710 460999 3712
rect 372889 3707 372955 3710
rect 460933 3707 460999 3710
rect 513281 3770 513347 3773
rect 516225 3770 516291 3773
rect 513281 3768 516291 3770
rect 513281 3712 513286 3768
rect 513342 3712 516230 3768
rect 516286 3712 516291 3768
rect 513281 3710 516291 3712
rect 513281 3707 513347 3710
rect 516225 3707 516291 3710
rect 518801 3770 518867 3773
rect 518985 3770 519051 3773
rect 518801 3768 519051 3770
rect 518801 3712 518806 3768
rect 518862 3712 518990 3768
rect 519046 3712 519051 3768
rect 518801 3710 519051 3712
rect 518801 3707 518867 3710
rect 518985 3707 519051 3710
rect 20621 3634 20687 3637
rect 161565 3634 161631 3637
rect 20621 3632 161631 3634
rect 20621 3576 20626 3632
rect 20682 3576 161570 3632
rect 161626 3576 161631 3632
rect 20621 3574 161631 3576
rect 20621 3571 20687 3574
rect 161565 3571 161631 3574
rect 369393 3634 369459 3637
rect 459645 3634 459711 3637
rect 369393 3632 459711 3634
rect 369393 3576 369398 3632
rect 369454 3576 459650 3632
rect 459706 3576 459711 3632
rect 369393 3574 459711 3576
rect 369393 3571 369459 3574
rect 459645 3571 459711 3574
rect 517421 3634 517487 3637
rect 582189 3634 582255 3637
rect 517421 3632 582255 3634
rect 517421 3576 517426 3632
rect 517482 3576 582194 3632
rect 582250 3576 582255 3632
rect 517421 3574 582255 3576
rect 517421 3571 517487 3574
rect 582189 3571 582255 3574
rect 11145 3498 11211 3501
rect 160277 3498 160343 3501
rect 11145 3496 160343 3498
rect 11145 3440 11150 3496
rect 11206 3440 160282 3496
rect 160338 3440 160343 3496
rect 11145 3438 160343 3440
rect 11145 3435 11211 3438
rect 160277 3435 160343 3438
rect 365805 3498 365871 3501
rect 459737 3498 459803 3501
rect 365805 3496 459803 3498
rect 365805 3440 365810 3496
rect 365866 3440 459742 3496
rect 459798 3440 459803 3496
rect 365805 3438 459803 3440
rect 365805 3435 365871 3438
rect 459737 3435 459803 3438
rect 514661 3498 514727 3501
rect 578601 3498 578667 3501
rect 514661 3496 578667 3498
rect 514661 3440 514666 3496
rect 514722 3440 578606 3496
rect 578662 3440 578667 3496
rect 514661 3438 578667 3440
rect 514661 3435 514727 3438
rect 578601 3435 578667 3438
rect 5257 3362 5323 3365
rect 164325 3362 164391 3365
rect 5257 3360 164391 3362
rect 5257 3304 5262 3360
rect 5318 3304 164330 3360
rect 164386 3304 164391 3360
rect 5257 3302 164391 3304
rect 5257 3299 5323 3302
rect 164325 3299 164391 3302
rect 362309 3362 362375 3365
rect 458173 3362 458239 3365
rect 362309 3360 458239 3362
rect 362309 3304 362314 3360
rect 362370 3304 458178 3360
rect 458234 3304 458239 3360
rect 362309 3302 458239 3304
rect 362309 3299 362375 3302
rect 458173 3299 458239 3302
rect 515857 3362 515923 3365
rect 580993 3362 581059 3365
rect 515857 3360 581059 3362
rect 515857 3304 515862 3360
rect 515918 3304 580998 3360
rect 581054 3304 581059 3360
rect 515857 3302 581059 3304
rect 515857 3299 515923 3302
rect 580993 3299 581059 3302
rect 460933 3090 460999 3093
rect 462313 3090 462379 3093
rect 460933 3088 462379 3090
rect 460933 3032 460938 3088
rect 460994 3032 462318 3088
rect 462374 3032 462379 3088
rect 460933 3030 462379 3032
rect 460933 3027 460999 3030
rect 462313 3027 462379 3030
rect 132217 2954 132283 2957
rect 134057 2954 134123 2957
rect 132217 2952 134123 2954
rect 132217 2896 132222 2952
rect 132278 2896 134062 2952
rect 134118 2896 134123 2952
rect 132217 2894 134123 2896
rect 132217 2891 132283 2894
rect 134057 2891 134123 2894
rect 128353 2818 128419 2821
rect 132585 2818 132651 2821
rect 128353 2816 132651 2818
rect 128353 2760 128358 2816
rect 128414 2760 132590 2816
rect 132646 2760 132651 2816
rect 128353 2758 132651 2760
rect 128353 2755 128419 2758
rect 132585 2755 132651 2758
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 12604 710478 13204 711440
rect 12604 710242 12786 710478
rect 13022 710242 13204 710478
rect 12604 710158 13204 710242
rect 12604 709922 12786 710158
rect 13022 709922 13204 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 9004 708598 9604 709560
rect 9004 708362 9186 708598
rect 9422 708362 9604 708598
rect 9004 708278 9604 708362
rect 9004 708042 9186 708278
rect 9422 708042 9604 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 5404 706718 6004 707680
rect 5404 706482 5586 706718
rect 5822 706482 6004 706718
rect 5404 706398 6004 706482
rect 5404 706162 5586 706398
rect 5822 706162 6004 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 699906 -2336 705222
rect -2936 699670 -2754 699906
rect -2518 699670 -2336 699906
rect -2936 699586 -2336 699670
rect -2936 699350 -2754 699586
rect -2518 699350 -2336 699586
rect -2936 684906 -2336 699350
rect -2936 684670 -2754 684906
rect -2518 684670 -2336 684906
rect -2936 684586 -2336 684670
rect -2936 684350 -2754 684586
rect -2518 684350 -2336 684586
rect -2936 669906 -2336 684350
rect -2936 669670 -2754 669906
rect -2518 669670 -2336 669906
rect -2936 669586 -2336 669670
rect -2936 669350 -2754 669586
rect -2518 669350 -2336 669586
rect -2936 -1286 -2336 669350
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 692406 -1396 704282
rect -1996 692170 -1814 692406
rect -1578 692170 -1396 692406
rect -1996 692086 -1396 692170
rect -1996 691850 -1814 692086
rect -1578 691850 -1396 692086
rect -1996 677406 -1396 691850
rect -1996 677170 -1814 677406
rect -1578 677170 -1396 677406
rect -1996 677086 -1396 677170
rect -1996 676850 -1814 677086
rect -1578 676850 -1396 677086
rect -1996 662406 -1396 676850
rect -1996 662170 -1814 662406
rect -1578 662170 -1396 662406
rect -1996 662086 -1396 662170
rect -1996 661850 -1814 662086
rect -1578 661850 -1396 662086
rect -1996 -346 -1396 661850
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 5404 -2226 6004 706162
rect 5404 -2462 5586 -2226
rect 5822 -2462 6004 -2226
rect 5404 -2546 6004 -2462
rect 5404 -2782 5586 -2546
rect 5822 -2782 6004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 5404 -3744 6004 -2782
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 9004 -4106 9604 708042
rect 9004 -4342 9186 -4106
rect 9422 -4342 9604 -4106
rect 9004 -4426 9604 -4342
rect 9004 -4662 9186 -4426
rect 9422 -4662 9604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 9004 -5624 9604 -4662
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 12604 -5986 13204 709922
rect 30604 711418 31204 711440
rect 30604 711182 30786 711418
rect 31022 711182 31204 711418
rect 30604 711098 31204 711182
rect 30604 710862 30786 711098
rect 31022 710862 31204 711098
rect 27004 709538 27604 709560
rect 27004 709302 27186 709538
rect 27422 709302 27604 709538
rect 27004 709218 27604 709302
rect 27004 708982 27186 709218
rect 27422 708982 27604 709218
rect 23404 707658 24004 707680
rect 23404 707422 23586 707658
rect 23822 707422 24004 707658
rect 23404 707338 24004 707422
rect 23404 707102 23586 707338
rect 23822 707102 24004 707338
rect 23404 -3166 24004 707102
rect 23404 -3402 23586 -3166
rect 23822 -3402 24004 -3166
rect 23404 -3486 24004 -3402
rect 23404 -3722 23586 -3486
rect 23822 -3722 24004 -3486
rect 23404 -3744 24004 -3722
rect 27004 -5046 27604 708982
rect 27004 -5282 27186 -5046
rect 27422 -5282 27604 -5046
rect 27004 -5366 27604 -5282
rect 27004 -5602 27186 -5366
rect 27422 -5602 27604 -5366
rect 27004 -5624 27604 -5602
rect 12604 -6222 12786 -5986
rect 13022 -6222 13204 -5986
rect 12604 -6306 13204 -6222
rect 12604 -6542 12786 -6306
rect 13022 -6542 13204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 12604 -7504 13204 -6542
rect 30604 -6926 31204 710862
rect 48604 710478 49204 711440
rect 48604 710242 48786 710478
rect 49022 710242 49204 710478
rect 48604 710158 49204 710242
rect 48604 709922 48786 710158
rect 49022 709922 49204 710158
rect 45004 708598 45604 709560
rect 45004 708362 45186 708598
rect 45422 708362 45604 708598
rect 45004 708278 45604 708362
rect 45004 708042 45186 708278
rect 45422 708042 45604 708278
rect 41404 706718 42004 707680
rect 41404 706482 41586 706718
rect 41822 706482 42004 706718
rect 41404 706398 42004 706482
rect 41404 706162 41586 706398
rect 41822 706162 42004 706398
rect 41404 -2226 42004 706162
rect 41404 -2462 41586 -2226
rect 41822 -2462 42004 -2226
rect 41404 -2546 42004 -2462
rect 41404 -2782 41586 -2546
rect 41822 -2782 42004 -2546
rect 41404 -3744 42004 -2782
rect 45004 -4106 45604 708042
rect 45004 -4342 45186 -4106
rect 45422 -4342 45604 -4106
rect 45004 -4426 45604 -4342
rect 45004 -4662 45186 -4426
rect 45422 -4662 45604 -4426
rect 45004 -5624 45604 -4662
rect 30604 -7162 30786 -6926
rect 31022 -7162 31204 -6926
rect 30604 -7246 31204 -7162
rect 30604 -7482 30786 -7246
rect 31022 -7482 31204 -7246
rect 30604 -7504 31204 -7482
rect 48604 -5986 49204 709922
rect 66604 711418 67204 711440
rect 66604 711182 66786 711418
rect 67022 711182 67204 711418
rect 66604 711098 67204 711182
rect 66604 710862 66786 711098
rect 67022 710862 67204 711098
rect 63004 709538 63604 709560
rect 63004 709302 63186 709538
rect 63422 709302 63604 709538
rect 63004 709218 63604 709302
rect 63004 708982 63186 709218
rect 63422 708982 63604 709218
rect 59404 707658 60004 707680
rect 59404 707422 59586 707658
rect 59822 707422 60004 707658
rect 59404 707338 60004 707422
rect 59404 707102 59586 707338
rect 59822 707102 60004 707338
rect 59404 -3166 60004 707102
rect 59404 -3402 59586 -3166
rect 59822 -3402 60004 -3166
rect 59404 -3486 60004 -3402
rect 59404 -3722 59586 -3486
rect 59822 -3722 60004 -3486
rect 59404 -3744 60004 -3722
rect 63004 -5046 63604 708982
rect 63004 -5282 63186 -5046
rect 63422 -5282 63604 -5046
rect 63004 -5366 63604 -5282
rect 63004 -5602 63186 -5366
rect 63422 -5602 63604 -5366
rect 63004 -5624 63604 -5602
rect 48604 -6222 48786 -5986
rect 49022 -6222 49204 -5986
rect 48604 -6306 49204 -6222
rect 48604 -6542 48786 -6306
rect 49022 -6542 49204 -6306
rect 48604 -7504 49204 -6542
rect 66604 -6926 67204 710862
rect 84604 710478 85204 711440
rect 84604 710242 84786 710478
rect 85022 710242 85204 710478
rect 84604 710158 85204 710242
rect 84604 709922 84786 710158
rect 85022 709922 85204 710158
rect 81004 708598 81604 709560
rect 81004 708362 81186 708598
rect 81422 708362 81604 708598
rect 81004 708278 81604 708362
rect 81004 708042 81186 708278
rect 81422 708042 81604 708278
rect 77404 706718 78004 707680
rect 77404 706482 77586 706718
rect 77822 706482 78004 706718
rect 77404 706398 78004 706482
rect 77404 706162 77586 706398
rect 77822 706162 78004 706398
rect 77404 682008 78004 706162
rect 81004 682008 81604 708042
rect 84604 682008 85204 709922
rect 102604 711418 103204 711440
rect 102604 711182 102786 711418
rect 103022 711182 103204 711418
rect 102604 711098 103204 711182
rect 102604 710862 102786 711098
rect 103022 710862 103204 711098
rect 99004 709538 99604 709560
rect 99004 709302 99186 709538
rect 99422 709302 99604 709538
rect 99004 709218 99604 709302
rect 99004 708982 99186 709218
rect 99422 708982 99604 709218
rect 95404 707658 96004 707680
rect 95404 707422 95586 707658
rect 95822 707422 96004 707658
rect 95404 707338 96004 707422
rect 95404 707102 95586 707338
rect 95822 707102 96004 707338
rect 95404 682008 96004 707102
rect 99004 682008 99604 708982
rect 102604 682008 103204 710862
rect 120604 710478 121204 711440
rect 120604 710242 120786 710478
rect 121022 710242 121204 710478
rect 120604 710158 121204 710242
rect 120604 709922 120786 710158
rect 121022 709922 121204 710158
rect 117004 708598 117604 709560
rect 117004 708362 117186 708598
rect 117422 708362 117604 708598
rect 117004 708278 117604 708362
rect 117004 708042 117186 708278
rect 117422 708042 117604 708278
rect 113404 706718 114004 707680
rect 113404 706482 113586 706718
rect 113822 706482 114004 706718
rect 113404 706398 114004 706482
rect 113404 706162 113586 706398
rect 113822 706162 114004 706398
rect 113404 682008 114004 706162
rect 117004 682008 117604 708042
rect 120604 682008 121204 709922
rect 138604 711418 139204 711440
rect 138604 711182 138786 711418
rect 139022 711182 139204 711418
rect 138604 711098 139204 711182
rect 138604 710862 138786 711098
rect 139022 710862 139204 711098
rect 135004 709538 135604 709560
rect 135004 709302 135186 709538
rect 135422 709302 135604 709538
rect 135004 709218 135604 709302
rect 135004 708982 135186 709218
rect 135422 708982 135604 709218
rect 131404 707658 132004 707680
rect 131404 707422 131586 707658
rect 131822 707422 132004 707658
rect 131404 707338 132004 707422
rect 131404 707102 131586 707338
rect 131822 707102 132004 707338
rect 131404 682008 132004 707102
rect 135004 682008 135604 708982
rect 138604 682008 139204 710862
rect 156604 710478 157204 711440
rect 156604 710242 156786 710478
rect 157022 710242 157204 710478
rect 156604 710158 157204 710242
rect 156604 709922 156786 710158
rect 157022 709922 157204 710158
rect 153004 708598 153604 709560
rect 153004 708362 153186 708598
rect 153422 708362 153604 708598
rect 153004 708278 153604 708362
rect 153004 708042 153186 708278
rect 153422 708042 153604 708278
rect 149404 706718 150004 707680
rect 149404 706482 149586 706718
rect 149822 706482 150004 706718
rect 149404 706398 150004 706482
rect 149404 706162 149586 706398
rect 149822 706162 150004 706398
rect 149404 682008 150004 706162
rect 153004 682008 153604 708042
rect 156604 682008 157204 709922
rect 174604 711418 175204 711440
rect 174604 711182 174786 711418
rect 175022 711182 175204 711418
rect 174604 711098 175204 711182
rect 174604 710862 174786 711098
rect 175022 710862 175204 711098
rect 171004 709538 171604 709560
rect 171004 709302 171186 709538
rect 171422 709302 171604 709538
rect 171004 709218 171604 709302
rect 171004 708982 171186 709218
rect 171422 708982 171604 709218
rect 167404 707658 168004 707680
rect 167404 707422 167586 707658
rect 167822 707422 168004 707658
rect 167404 707338 168004 707422
rect 167404 707102 167586 707338
rect 167822 707102 168004 707338
rect 167404 682008 168004 707102
rect 171004 682008 171604 708982
rect 174604 682008 175204 710862
rect 192604 710478 193204 711440
rect 192604 710242 192786 710478
rect 193022 710242 193204 710478
rect 192604 710158 193204 710242
rect 192604 709922 192786 710158
rect 193022 709922 193204 710158
rect 189004 708598 189604 709560
rect 189004 708362 189186 708598
rect 189422 708362 189604 708598
rect 189004 708278 189604 708362
rect 189004 708042 189186 708278
rect 189422 708042 189604 708278
rect 185404 706718 186004 707680
rect 185404 706482 185586 706718
rect 185822 706482 186004 706718
rect 185404 706398 186004 706482
rect 185404 706162 185586 706398
rect 185822 706162 186004 706398
rect 185404 682008 186004 706162
rect 189004 682008 189604 708042
rect 192604 682008 193204 709922
rect 210604 711418 211204 711440
rect 210604 711182 210786 711418
rect 211022 711182 211204 711418
rect 210604 711098 211204 711182
rect 210604 710862 210786 711098
rect 211022 710862 211204 711098
rect 207004 709538 207604 709560
rect 207004 709302 207186 709538
rect 207422 709302 207604 709538
rect 207004 709218 207604 709302
rect 207004 708982 207186 709218
rect 207422 708982 207604 709218
rect 203404 707658 204004 707680
rect 203404 707422 203586 707658
rect 203822 707422 204004 707658
rect 203404 707338 204004 707422
rect 203404 707102 203586 707338
rect 203822 707102 204004 707338
rect 203404 682008 204004 707102
rect 207004 682008 207604 708982
rect 210604 682008 211204 710862
rect 228604 710478 229204 711440
rect 228604 710242 228786 710478
rect 229022 710242 229204 710478
rect 228604 710158 229204 710242
rect 228604 709922 228786 710158
rect 229022 709922 229204 710158
rect 225004 708598 225604 709560
rect 225004 708362 225186 708598
rect 225422 708362 225604 708598
rect 225004 708278 225604 708362
rect 225004 708042 225186 708278
rect 225422 708042 225604 708278
rect 221404 706718 222004 707680
rect 221404 706482 221586 706718
rect 221822 706482 222004 706718
rect 221404 706398 222004 706482
rect 221404 706162 221586 706398
rect 221822 706162 222004 706398
rect 221404 682008 222004 706162
rect 225004 682008 225604 708042
rect 228604 682008 229204 709922
rect 246604 711418 247204 711440
rect 246604 711182 246786 711418
rect 247022 711182 247204 711418
rect 246604 711098 247204 711182
rect 246604 710862 246786 711098
rect 247022 710862 247204 711098
rect 243004 709538 243604 709560
rect 243004 709302 243186 709538
rect 243422 709302 243604 709538
rect 243004 709218 243604 709302
rect 243004 708982 243186 709218
rect 243422 708982 243604 709218
rect 239404 707658 240004 707680
rect 239404 707422 239586 707658
rect 239822 707422 240004 707658
rect 239404 707338 240004 707422
rect 239404 707102 239586 707338
rect 239822 707102 240004 707338
rect 239404 682008 240004 707102
rect 243004 682008 243604 708982
rect 246604 682008 247204 710862
rect 264604 710478 265204 711440
rect 264604 710242 264786 710478
rect 265022 710242 265204 710478
rect 264604 710158 265204 710242
rect 264604 709922 264786 710158
rect 265022 709922 265204 710158
rect 261004 708598 261604 709560
rect 261004 708362 261186 708598
rect 261422 708362 261604 708598
rect 261004 708278 261604 708362
rect 261004 708042 261186 708278
rect 261422 708042 261604 708278
rect 257404 706718 258004 707680
rect 257404 706482 257586 706718
rect 257822 706482 258004 706718
rect 257404 706398 258004 706482
rect 257404 706162 257586 706398
rect 257822 706162 258004 706398
rect 257404 682008 258004 706162
rect 261004 682008 261604 708042
rect 264604 682008 265204 709922
rect 282604 711418 283204 711440
rect 282604 711182 282786 711418
rect 283022 711182 283204 711418
rect 282604 711098 283204 711182
rect 282604 710862 282786 711098
rect 283022 710862 283204 711098
rect 279004 709538 279604 709560
rect 279004 709302 279186 709538
rect 279422 709302 279604 709538
rect 279004 709218 279604 709302
rect 279004 708982 279186 709218
rect 279422 708982 279604 709218
rect 275404 707658 276004 707680
rect 275404 707422 275586 707658
rect 275822 707422 276004 707658
rect 275404 707338 276004 707422
rect 275404 707102 275586 707338
rect 275822 707102 276004 707338
rect 275404 682008 276004 707102
rect 279004 682008 279604 708982
rect 282604 682008 283204 710862
rect 300604 710478 301204 711440
rect 300604 710242 300786 710478
rect 301022 710242 301204 710478
rect 300604 710158 301204 710242
rect 300604 709922 300786 710158
rect 301022 709922 301204 710158
rect 297004 708598 297604 709560
rect 297004 708362 297186 708598
rect 297422 708362 297604 708598
rect 297004 708278 297604 708362
rect 297004 708042 297186 708278
rect 297422 708042 297604 708278
rect 293404 706718 294004 707680
rect 293404 706482 293586 706718
rect 293822 706482 294004 706718
rect 293404 706398 294004 706482
rect 293404 706162 293586 706398
rect 293822 706162 294004 706398
rect 293404 682008 294004 706162
rect 297004 682008 297604 708042
rect 300604 682008 301204 709922
rect 318604 711418 319204 711440
rect 318604 711182 318786 711418
rect 319022 711182 319204 711418
rect 318604 711098 319204 711182
rect 318604 710862 318786 711098
rect 319022 710862 319204 711098
rect 315004 709538 315604 709560
rect 315004 709302 315186 709538
rect 315422 709302 315604 709538
rect 315004 709218 315604 709302
rect 315004 708982 315186 709218
rect 315422 708982 315604 709218
rect 311404 707658 312004 707680
rect 311404 707422 311586 707658
rect 311822 707422 312004 707658
rect 311404 707338 312004 707422
rect 311404 707102 311586 707338
rect 311822 707102 312004 707338
rect 311404 682008 312004 707102
rect 315004 682008 315604 708982
rect 318604 682008 319204 710862
rect 336604 710478 337204 711440
rect 336604 710242 336786 710478
rect 337022 710242 337204 710478
rect 336604 710158 337204 710242
rect 336604 709922 336786 710158
rect 337022 709922 337204 710158
rect 333004 708598 333604 709560
rect 333004 708362 333186 708598
rect 333422 708362 333604 708598
rect 333004 708278 333604 708362
rect 333004 708042 333186 708278
rect 333422 708042 333604 708278
rect 329404 706718 330004 707680
rect 329404 706482 329586 706718
rect 329822 706482 330004 706718
rect 329404 706398 330004 706482
rect 329404 706162 329586 706398
rect 329822 706162 330004 706398
rect 329404 682008 330004 706162
rect 333004 682008 333604 708042
rect 336604 682008 337204 709922
rect 354604 711418 355204 711440
rect 354604 711182 354786 711418
rect 355022 711182 355204 711418
rect 354604 711098 355204 711182
rect 354604 710862 354786 711098
rect 355022 710862 355204 711098
rect 351004 709538 351604 709560
rect 351004 709302 351186 709538
rect 351422 709302 351604 709538
rect 351004 709218 351604 709302
rect 351004 708982 351186 709218
rect 351422 708982 351604 709218
rect 347404 707658 348004 707680
rect 347404 707422 347586 707658
rect 347822 707422 348004 707658
rect 347404 707338 348004 707422
rect 347404 707102 347586 707338
rect 347822 707102 348004 707338
rect 347404 682008 348004 707102
rect 351004 682008 351604 708982
rect 354604 682008 355204 710862
rect 372604 710478 373204 711440
rect 372604 710242 372786 710478
rect 373022 710242 373204 710478
rect 372604 710158 373204 710242
rect 372604 709922 372786 710158
rect 373022 709922 373204 710158
rect 369004 708598 369604 709560
rect 369004 708362 369186 708598
rect 369422 708362 369604 708598
rect 369004 708278 369604 708362
rect 369004 708042 369186 708278
rect 369422 708042 369604 708278
rect 365404 706718 366004 707680
rect 365404 706482 365586 706718
rect 365822 706482 366004 706718
rect 365404 706398 366004 706482
rect 365404 706162 365586 706398
rect 365822 706162 366004 706398
rect 365404 682008 366004 706162
rect 369004 682008 369604 708042
rect 372604 682008 373204 709922
rect 390604 711418 391204 711440
rect 390604 711182 390786 711418
rect 391022 711182 391204 711418
rect 390604 711098 391204 711182
rect 390604 710862 390786 711098
rect 391022 710862 391204 711098
rect 387004 709538 387604 709560
rect 387004 709302 387186 709538
rect 387422 709302 387604 709538
rect 387004 709218 387604 709302
rect 387004 708982 387186 709218
rect 387422 708982 387604 709218
rect 383404 707658 384004 707680
rect 383404 707422 383586 707658
rect 383822 707422 384004 707658
rect 383404 707338 384004 707422
rect 383404 707102 383586 707338
rect 383822 707102 384004 707338
rect 383404 682008 384004 707102
rect 387004 682008 387604 708982
rect 390604 682008 391204 710862
rect 408604 710478 409204 711440
rect 408604 710242 408786 710478
rect 409022 710242 409204 710478
rect 408604 710158 409204 710242
rect 408604 709922 408786 710158
rect 409022 709922 409204 710158
rect 405004 708598 405604 709560
rect 405004 708362 405186 708598
rect 405422 708362 405604 708598
rect 405004 708278 405604 708362
rect 405004 708042 405186 708278
rect 405422 708042 405604 708278
rect 401404 706718 402004 707680
rect 401404 706482 401586 706718
rect 401822 706482 402004 706718
rect 401404 706398 402004 706482
rect 401404 706162 401586 706398
rect 401822 706162 402004 706398
rect 401404 682008 402004 706162
rect 405004 682008 405604 708042
rect 408604 682008 409204 709922
rect 426604 711418 427204 711440
rect 426604 711182 426786 711418
rect 427022 711182 427204 711418
rect 426604 711098 427204 711182
rect 426604 710862 426786 711098
rect 427022 710862 427204 711098
rect 423004 709538 423604 709560
rect 423004 709302 423186 709538
rect 423422 709302 423604 709538
rect 423004 709218 423604 709302
rect 423004 708982 423186 709218
rect 423422 708982 423604 709218
rect 419404 707658 420004 707680
rect 419404 707422 419586 707658
rect 419822 707422 420004 707658
rect 419404 707338 420004 707422
rect 419404 707102 419586 707338
rect 419822 707102 420004 707338
rect 419404 682008 420004 707102
rect 423004 682008 423604 708982
rect 426604 682008 427204 710862
rect 444604 710478 445204 711440
rect 444604 710242 444786 710478
rect 445022 710242 445204 710478
rect 444604 710158 445204 710242
rect 444604 709922 444786 710158
rect 445022 709922 445204 710158
rect 441004 708598 441604 709560
rect 441004 708362 441186 708598
rect 441422 708362 441604 708598
rect 441004 708278 441604 708362
rect 441004 708042 441186 708278
rect 441422 708042 441604 708278
rect 437404 706718 438004 707680
rect 437404 706482 437586 706718
rect 437822 706482 438004 706718
rect 437404 706398 438004 706482
rect 437404 706162 437586 706398
rect 437822 706162 438004 706398
rect 437404 682008 438004 706162
rect 441004 682008 441604 708042
rect 444604 682008 445204 709922
rect 462604 711418 463204 711440
rect 462604 711182 462786 711418
rect 463022 711182 463204 711418
rect 462604 711098 463204 711182
rect 462604 710862 462786 711098
rect 463022 710862 463204 711098
rect 459004 709538 459604 709560
rect 459004 709302 459186 709538
rect 459422 709302 459604 709538
rect 459004 709218 459604 709302
rect 459004 708982 459186 709218
rect 459422 708982 459604 709218
rect 455404 707658 456004 707680
rect 455404 707422 455586 707658
rect 455822 707422 456004 707658
rect 455404 707338 456004 707422
rect 455404 707102 455586 707338
rect 455822 707102 456004 707338
rect 455404 682008 456004 707102
rect 459004 682008 459604 708982
rect 462604 682008 463204 710862
rect 480604 710478 481204 711440
rect 480604 710242 480786 710478
rect 481022 710242 481204 710478
rect 480604 710158 481204 710242
rect 480604 709922 480786 710158
rect 481022 709922 481204 710158
rect 477004 708598 477604 709560
rect 477004 708362 477186 708598
rect 477422 708362 477604 708598
rect 477004 708278 477604 708362
rect 477004 708042 477186 708278
rect 477422 708042 477604 708278
rect 473404 706718 474004 707680
rect 473404 706482 473586 706718
rect 473822 706482 474004 706718
rect 473404 706398 474004 706482
rect 473404 706162 473586 706398
rect 473822 706162 474004 706398
rect 473404 682008 474004 706162
rect 477004 682008 477604 708042
rect 480604 682008 481204 709922
rect 498604 711418 499204 711440
rect 498604 711182 498786 711418
rect 499022 711182 499204 711418
rect 498604 711098 499204 711182
rect 498604 710862 498786 711098
rect 499022 710862 499204 711098
rect 495004 709538 495604 709560
rect 495004 709302 495186 709538
rect 495422 709302 495604 709538
rect 495004 709218 495604 709302
rect 495004 708982 495186 709218
rect 495422 708982 495604 709218
rect 491404 707658 492004 707680
rect 491404 707422 491586 707658
rect 491822 707422 492004 707658
rect 491404 707338 492004 707422
rect 491404 707102 491586 707338
rect 491822 707102 492004 707338
rect 491404 682008 492004 707102
rect 495004 682008 495604 708982
rect 498604 682008 499204 710862
rect 516604 710478 517204 711440
rect 516604 710242 516786 710478
rect 517022 710242 517204 710478
rect 516604 710158 517204 710242
rect 516604 709922 516786 710158
rect 517022 709922 517204 710158
rect 513004 708598 513604 709560
rect 513004 708362 513186 708598
rect 513422 708362 513604 708598
rect 513004 708278 513604 708362
rect 513004 708042 513186 708278
rect 513422 708042 513604 708278
rect 509404 706718 510004 707680
rect 509404 706482 509586 706718
rect 509822 706482 510004 706718
rect 509404 706398 510004 706482
rect 509404 706162 509586 706398
rect 509822 706162 510004 706398
rect 509404 682008 510004 706162
rect 513004 682008 513604 708042
rect 516604 682008 517204 709922
rect 534604 711418 535204 711440
rect 534604 711182 534786 711418
rect 535022 711182 535204 711418
rect 534604 711098 535204 711182
rect 534604 710862 534786 711098
rect 535022 710862 535204 711098
rect 531004 709538 531604 709560
rect 531004 709302 531186 709538
rect 531422 709302 531604 709538
rect 531004 709218 531604 709302
rect 531004 708982 531186 709218
rect 531422 708982 531604 709218
rect 527404 707658 528004 707680
rect 527404 707422 527586 707658
rect 527822 707422 528004 707658
rect 527404 707338 528004 707422
rect 527404 707102 527586 707338
rect 527822 707102 528004 707338
rect 72158 677406 72958 677428
rect 72158 677170 72280 677406
rect 72516 677170 72600 677406
rect 72836 677170 72958 677406
rect 72158 677086 72958 677170
rect 72158 676850 72280 677086
rect 72516 676850 72600 677086
rect 72836 676850 72958 677086
rect 72158 676828 72958 676850
rect 514990 677406 515790 677428
rect 514990 677170 515112 677406
rect 515348 677170 515432 677406
rect 515668 677170 515790 677406
rect 514990 677086 515790 677170
rect 514990 676850 515112 677086
rect 515348 676850 515432 677086
rect 515668 676850 515790 677086
rect 514990 676828 515790 676850
rect 70998 669906 71798 669928
rect 70998 669670 71120 669906
rect 71356 669670 71440 669906
rect 71676 669670 71798 669906
rect 70998 669586 71798 669670
rect 70998 669350 71120 669586
rect 71356 669350 71440 669586
rect 71676 669350 71798 669586
rect 70998 669328 71798 669350
rect 516150 669906 516950 669928
rect 516150 669670 516272 669906
rect 516508 669670 516592 669906
rect 516828 669670 516950 669906
rect 516150 669586 516950 669670
rect 516150 669350 516272 669586
rect 516508 669350 516592 669586
rect 516828 669350 516950 669586
rect 516150 669328 516950 669350
rect 72158 662406 72958 662428
rect 72158 662170 72280 662406
rect 72516 662170 72600 662406
rect 72836 662170 72958 662406
rect 72158 662086 72958 662170
rect 72158 661850 72280 662086
rect 72516 661850 72600 662086
rect 72836 661850 72958 662086
rect 72158 661828 72958 661850
rect 514990 662406 515790 662428
rect 514990 662170 515112 662406
rect 515348 662170 515432 662406
rect 515668 662170 515790 662406
rect 514990 662086 515790 662170
rect 514990 661850 515112 662086
rect 515348 661850 515432 662086
rect 515668 661850 515790 662086
rect 514990 661828 515790 661850
rect 77404 -2226 78004 86000
rect 77404 -2462 77586 -2226
rect 77822 -2462 78004 -2226
rect 77404 -2546 78004 -2462
rect 77404 -2782 77586 -2546
rect 77822 -2782 78004 -2546
rect 77404 -3744 78004 -2782
rect 81004 -4106 81604 86000
rect 81004 -4342 81186 -4106
rect 81422 -4342 81604 -4106
rect 81004 -4426 81604 -4342
rect 81004 -4662 81186 -4426
rect 81422 -4662 81604 -4426
rect 81004 -5624 81604 -4662
rect 66604 -7162 66786 -6926
rect 67022 -7162 67204 -6926
rect 66604 -7246 67204 -7162
rect 66604 -7482 66786 -7246
rect 67022 -7482 67204 -7246
rect 66604 -7504 67204 -7482
rect 84604 -5986 85204 86000
rect 95404 -3166 96004 86000
rect 95404 -3402 95586 -3166
rect 95822 -3402 96004 -3166
rect 95404 -3486 96004 -3402
rect 95404 -3722 95586 -3486
rect 95822 -3722 96004 -3486
rect 95404 -3744 96004 -3722
rect 99004 -5046 99604 86000
rect 99004 -5282 99186 -5046
rect 99422 -5282 99604 -5046
rect 99004 -5366 99604 -5282
rect 99004 -5602 99186 -5366
rect 99422 -5602 99604 -5366
rect 99004 -5624 99604 -5602
rect 84604 -6222 84786 -5986
rect 85022 -6222 85204 -5986
rect 84604 -6306 85204 -6222
rect 84604 -6542 84786 -6306
rect 85022 -6542 85204 -6306
rect 84604 -7504 85204 -6542
rect 102604 -6926 103204 86000
rect 113404 -2226 114004 86000
rect 113404 -2462 113586 -2226
rect 113822 -2462 114004 -2226
rect 113404 -2546 114004 -2462
rect 113404 -2782 113586 -2546
rect 113822 -2782 114004 -2546
rect 113404 -3744 114004 -2782
rect 117004 -4106 117604 86000
rect 117004 -4342 117186 -4106
rect 117422 -4342 117604 -4106
rect 117004 -4426 117604 -4342
rect 117004 -4662 117186 -4426
rect 117422 -4662 117604 -4426
rect 117004 -5624 117604 -4662
rect 102604 -7162 102786 -6926
rect 103022 -7162 103204 -6926
rect 102604 -7246 103204 -7162
rect 102604 -7482 102786 -7246
rect 103022 -7482 103204 -7246
rect 102604 -7504 103204 -7482
rect 120604 -5986 121204 86000
rect 131404 -3166 132004 86000
rect 131404 -3402 131586 -3166
rect 131822 -3402 132004 -3166
rect 131404 -3486 132004 -3402
rect 131404 -3722 131586 -3486
rect 131822 -3722 132004 -3486
rect 131404 -3744 132004 -3722
rect 135004 -5046 135604 86000
rect 135004 -5282 135186 -5046
rect 135422 -5282 135604 -5046
rect 135004 -5366 135604 -5282
rect 135004 -5602 135186 -5366
rect 135422 -5602 135604 -5366
rect 135004 -5624 135604 -5602
rect 120604 -6222 120786 -5986
rect 121022 -6222 121204 -5986
rect 120604 -6306 121204 -6222
rect 120604 -6542 120786 -6306
rect 121022 -6542 121204 -6306
rect 120604 -7504 121204 -6542
rect 138604 -6926 139204 86000
rect 149404 -2226 150004 86000
rect 149404 -2462 149586 -2226
rect 149822 -2462 150004 -2226
rect 149404 -2546 150004 -2462
rect 149404 -2782 149586 -2546
rect 149822 -2782 150004 -2546
rect 149404 -3744 150004 -2782
rect 153004 -4106 153604 86000
rect 153004 -4342 153186 -4106
rect 153422 -4342 153604 -4106
rect 153004 -4426 153604 -4342
rect 153004 -4662 153186 -4426
rect 153422 -4662 153604 -4426
rect 153004 -5624 153604 -4662
rect 138604 -7162 138786 -6926
rect 139022 -7162 139204 -6926
rect 138604 -7246 139204 -7162
rect 138604 -7482 138786 -7246
rect 139022 -7482 139204 -7246
rect 138604 -7504 139204 -7482
rect 156604 -5986 157204 86000
rect 167404 -3166 168004 86000
rect 167404 -3402 167586 -3166
rect 167822 -3402 168004 -3166
rect 167404 -3486 168004 -3402
rect 167404 -3722 167586 -3486
rect 167822 -3722 168004 -3486
rect 167404 -3744 168004 -3722
rect 171004 -5046 171604 86000
rect 171004 -5282 171186 -5046
rect 171422 -5282 171604 -5046
rect 171004 -5366 171604 -5282
rect 171004 -5602 171186 -5366
rect 171422 -5602 171604 -5366
rect 171004 -5624 171604 -5602
rect 156604 -6222 156786 -5986
rect 157022 -6222 157204 -5986
rect 156604 -6306 157204 -6222
rect 156604 -6542 156786 -6306
rect 157022 -6542 157204 -6306
rect 156604 -7504 157204 -6542
rect 174604 -6926 175204 86000
rect 185404 -2226 186004 86000
rect 185404 -2462 185586 -2226
rect 185822 -2462 186004 -2226
rect 185404 -2546 186004 -2462
rect 185404 -2782 185586 -2546
rect 185822 -2782 186004 -2546
rect 185404 -3744 186004 -2782
rect 189004 -4106 189604 86000
rect 189004 -4342 189186 -4106
rect 189422 -4342 189604 -4106
rect 189004 -4426 189604 -4342
rect 189004 -4662 189186 -4426
rect 189422 -4662 189604 -4426
rect 189004 -5624 189604 -4662
rect 174604 -7162 174786 -6926
rect 175022 -7162 175204 -6926
rect 174604 -7246 175204 -7162
rect 174604 -7482 174786 -7246
rect 175022 -7482 175204 -7246
rect 174604 -7504 175204 -7482
rect 192604 -5986 193204 86000
rect 203404 -3166 204004 86000
rect 203404 -3402 203586 -3166
rect 203822 -3402 204004 -3166
rect 203404 -3486 204004 -3402
rect 203404 -3722 203586 -3486
rect 203822 -3722 204004 -3486
rect 203404 -3744 204004 -3722
rect 207004 -5046 207604 86000
rect 207004 -5282 207186 -5046
rect 207422 -5282 207604 -5046
rect 207004 -5366 207604 -5282
rect 207004 -5602 207186 -5366
rect 207422 -5602 207604 -5366
rect 207004 -5624 207604 -5602
rect 192604 -6222 192786 -5986
rect 193022 -6222 193204 -5986
rect 192604 -6306 193204 -6222
rect 192604 -6542 192786 -6306
rect 193022 -6542 193204 -6306
rect 192604 -7504 193204 -6542
rect 210604 -6926 211204 86000
rect 221404 -2226 222004 86000
rect 221404 -2462 221586 -2226
rect 221822 -2462 222004 -2226
rect 221404 -2546 222004 -2462
rect 221404 -2782 221586 -2546
rect 221822 -2782 222004 -2546
rect 221404 -3744 222004 -2782
rect 225004 -4106 225604 86000
rect 225004 -4342 225186 -4106
rect 225422 -4342 225604 -4106
rect 225004 -4426 225604 -4342
rect 225004 -4662 225186 -4426
rect 225422 -4662 225604 -4426
rect 225004 -5624 225604 -4662
rect 210604 -7162 210786 -6926
rect 211022 -7162 211204 -6926
rect 210604 -7246 211204 -7162
rect 210604 -7482 210786 -7246
rect 211022 -7482 211204 -7246
rect 210604 -7504 211204 -7482
rect 228604 -5986 229204 86000
rect 239404 -3166 240004 86000
rect 239404 -3402 239586 -3166
rect 239822 -3402 240004 -3166
rect 239404 -3486 240004 -3402
rect 239404 -3722 239586 -3486
rect 239822 -3722 240004 -3486
rect 239404 -3744 240004 -3722
rect 243004 -5046 243604 86000
rect 243004 -5282 243186 -5046
rect 243422 -5282 243604 -5046
rect 243004 -5366 243604 -5282
rect 243004 -5602 243186 -5366
rect 243422 -5602 243604 -5366
rect 243004 -5624 243604 -5602
rect 228604 -6222 228786 -5986
rect 229022 -6222 229204 -5986
rect 228604 -6306 229204 -6222
rect 228604 -6542 228786 -6306
rect 229022 -6542 229204 -6306
rect 228604 -7504 229204 -6542
rect 246604 -6926 247204 86000
rect 257404 -2226 258004 86000
rect 257404 -2462 257586 -2226
rect 257822 -2462 258004 -2226
rect 257404 -2546 258004 -2462
rect 257404 -2782 257586 -2546
rect 257822 -2782 258004 -2546
rect 257404 -3744 258004 -2782
rect 261004 -4106 261604 86000
rect 261004 -4342 261186 -4106
rect 261422 -4342 261604 -4106
rect 261004 -4426 261604 -4342
rect 261004 -4662 261186 -4426
rect 261422 -4662 261604 -4426
rect 261004 -5624 261604 -4662
rect 246604 -7162 246786 -6926
rect 247022 -7162 247204 -6926
rect 246604 -7246 247204 -7162
rect 246604 -7482 246786 -7246
rect 247022 -7482 247204 -7246
rect 246604 -7504 247204 -7482
rect 264604 -5986 265204 86000
rect 275404 -3166 276004 86000
rect 275404 -3402 275586 -3166
rect 275822 -3402 276004 -3166
rect 275404 -3486 276004 -3402
rect 275404 -3722 275586 -3486
rect 275822 -3722 276004 -3486
rect 275404 -3744 276004 -3722
rect 279004 -5046 279604 86000
rect 279004 -5282 279186 -5046
rect 279422 -5282 279604 -5046
rect 279004 -5366 279604 -5282
rect 279004 -5602 279186 -5366
rect 279422 -5602 279604 -5366
rect 279004 -5624 279604 -5602
rect 264604 -6222 264786 -5986
rect 265022 -6222 265204 -5986
rect 264604 -6306 265204 -6222
rect 264604 -6542 264786 -6306
rect 265022 -6542 265204 -6306
rect 264604 -7504 265204 -6542
rect 282604 -6926 283204 86000
rect 293404 -2226 294004 86000
rect 293404 -2462 293586 -2226
rect 293822 -2462 294004 -2226
rect 293404 -2546 294004 -2462
rect 293404 -2782 293586 -2546
rect 293822 -2782 294004 -2546
rect 293404 -3744 294004 -2782
rect 297004 -4106 297604 86000
rect 297004 -4342 297186 -4106
rect 297422 -4342 297604 -4106
rect 297004 -4426 297604 -4342
rect 297004 -4662 297186 -4426
rect 297422 -4662 297604 -4426
rect 297004 -5624 297604 -4662
rect 282604 -7162 282786 -6926
rect 283022 -7162 283204 -6926
rect 282604 -7246 283204 -7162
rect 282604 -7482 282786 -7246
rect 283022 -7482 283204 -7246
rect 282604 -7504 283204 -7482
rect 300604 -5986 301204 86000
rect 311404 -3166 312004 86000
rect 311404 -3402 311586 -3166
rect 311822 -3402 312004 -3166
rect 311404 -3486 312004 -3402
rect 311404 -3722 311586 -3486
rect 311822 -3722 312004 -3486
rect 311404 -3744 312004 -3722
rect 315004 -5046 315604 86000
rect 315004 -5282 315186 -5046
rect 315422 -5282 315604 -5046
rect 315004 -5366 315604 -5282
rect 315004 -5602 315186 -5366
rect 315422 -5602 315604 -5366
rect 315004 -5624 315604 -5602
rect 300604 -6222 300786 -5986
rect 301022 -6222 301204 -5986
rect 300604 -6306 301204 -6222
rect 300604 -6542 300786 -6306
rect 301022 -6542 301204 -6306
rect 300604 -7504 301204 -6542
rect 318604 -6926 319204 86000
rect 329404 -2226 330004 86000
rect 329404 -2462 329586 -2226
rect 329822 -2462 330004 -2226
rect 329404 -2546 330004 -2462
rect 329404 -2782 329586 -2546
rect 329822 -2782 330004 -2546
rect 329404 -3744 330004 -2782
rect 333004 -4106 333604 86000
rect 333004 -4342 333186 -4106
rect 333422 -4342 333604 -4106
rect 333004 -4426 333604 -4342
rect 333004 -4662 333186 -4426
rect 333422 -4662 333604 -4426
rect 333004 -5624 333604 -4662
rect 318604 -7162 318786 -6926
rect 319022 -7162 319204 -6926
rect 318604 -7246 319204 -7162
rect 318604 -7482 318786 -7246
rect 319022 -7482 319204 -7246
rect 318604 -7504 319204 -7482
rect 336604 -5986 337204 86000
rect 347404 -3166 348004 86000
rect 347404 -3402 347586 -3166
rect 347822 -3402 348004 -3166
rect 347404 -3486 348004 -3402
rect 347404 -3722 347586 -3486
rect 347822 -3722 348004 -3486
rect 347404 -3744 348004 -3722
rect 351004 -5046 351604 86000
rect 351004 -5282 351186 -5046
rect 351422 -5282 351604 -5046
rect 351004 -5366 351604 -5282
rect 351004 -5602 351186 -5366
rect 351422 -5602 351604 -5366
rect 351004 -5624 351604 -5602
rect 336604 -6222 336786 -5986
rect 337022 -6222 337204 -5986
rect 336604 -6306 337204 -6222
rect 336604 -6542 336786 -6306
rect 337022 -6542 337204 -6306
rect 336604 -7504 337204 -6542
rect 354604 -6926 355204 86000
rect 365404 -2226 366004 86000
rect 365404 -2462 365586 -2226
rect 365822 -2462 366004 -2226
rect 365404 -2546 366004 -2462
rect 365404 -2782 365586 -2546
rect 365822 -2782 366004 -2546
rect 365404 -3744 366004 -2782
rect 369004 -4106 369604 86000
rect 369004 -4342 369186 -4106
rect 369422 -4342 369604 -4106
rect 369004 -4426 369604 -4342
rect 369004 -4662 369186 -4426
rect 369422 -4662 369604 -4426
rect 369004 -5624 369604 -4662
rect 354604 -7162 354786 -6926
rect 355022 -7162 355204 -6926
rect 354604 -7246 355204 -7162
rect 354604 -7482 354786 -7246
rect 355022 -7482 355204 -7246
rect 354604 -7504 355204 -7482
rect 372604 -5986 373204 86000
rect 383404 -3166 384004 86000
rect 383404 -3402 383586 -3166
rect 383822 -3402 384004 -3166
rect 383404 -3486 384004 -3402
rect 383404 -3722 383586 -3486
rect 383822 -3722 384004 -3486
rect 383404 -3744 384004 -3722
rect 387004 -5046 387604 86000
rect 387004 -5282 387186 -5046
rect 387422 -5282 387604 -5046
rect 387004 -5366 387604 -5282
rect 387004 -5602 387186 -5366
rect 387422 -5602 387604 -5366
rect 387004 -5624 387604 -5602
rect 372604 -6222 372786 -5986
rect 373022 -6222 373204 -5986
rect 372604 -6306 373204 -6222
rect 372604 -6542 372786 -6306
rect 373022 -6542 373204 -6306
rect 372604 -7504 373204 -6542
rect 390604 -6926 391204 86000
rect 401404 -2226 402004 86000
rect 401404 -2462 401586 -2226
rect 401822 -2462 402004 -2226
rect 401404 -2546 402004 -2462
rect 401404 -2782 401586 -2546
rect 401822 -2782 402004 -2546
rect 401404 -3744 402004 -2782
rect 405004 -4106 405604 86000
rect 405004 -4342 405186 -4106
rect 405422 -4342 405604 -4106
rect 405004 -4426 405604 -4342
rect 405004 -4662 405186 -4426
rect 405422 -4662 405604 -4426
rect 405004 -5624 405604 -4662
rect 390604 -7162 390786 -6926
rect 391022 -7162 391204 -6926
rect 390604 -7246 391204 -7162
rect 390604 -7482 390786 -7246
rect 391022 -7482 391204 -7246
rect 390604 -7504 391204 -7482
rect 408604 -5986 409204 86000
rect 419404 -3166 420004 86000
rect 419404 -3402 419586 -3166
rect 419822 -3402 420004 -3166
rect 419404 -3486 420004 -3402
rect 419404 -3722 419586 -3486
rect 419822 -3722 420004 -3486
rect 419404 -3744 420004 -3722
rect 423004 -5046 423604 86000
rect 423004 -5282 423186 -5046
rect 423422 -5282 423604 -5046
rect 423004 -5366 423604 -5282
rect 423004 -5602 423186 -5366
rect 423422 -5602 423604 -5366
rect 423004 -5624 423604 -5602
rect 408604 -6222 408786 -5986
rect 409022 -6222 409204 -5986
rect 408604 -6306 409204 -6222
rect 408604 -6542 408786 -6306
rect 409022 -6542 409204 -6306
rect 408604 -7504 409204 -6542
rect 426604 -6926 427204 86000
rect 437404 -2226 438004 86000
rect 437404 -2462 437586 -2226
rect 437822 -2462 438004 -2226
rect 437404 -2546 438004 -2462
rect 437404 -2782 437586 -2546
rect 437822 -2782 438004 -2546
rect 437404 -3744 438004 -2782
rect 441004 -4106 441604 86000
rect 441004 -4342 441186 -4106
rect 441422 -4342 441604 -4106
rect 441004 -4426 441604 -4342
rect 441004 -4662 441186 -4426
rect 441422 -4662 441604 -4426
rect 441004 -5624 441604 -4662
rect 426604 -7162 426786 -6926
rect 427022 -7162 427204 -6926
rect 426604 -7246 427204 -7162
rect 426604 -7482 426786 -7246
rect 427022 -7482 427204 -7246
rect 426604 -7504 427204 -7482
rect 444604 -5986 445204 86000
rect 455404 -3166 456004 86000
rect 455404 -3402 455586 -3166
rect 455822 -3402 456004 -3166
rect 455404 -3486 456004 -3402
rect 455404 -3722 455586 -3486
rect 455822 -3722 456004 -3486
rect 455404 -3744 456004 -3722
rect 459004 -5046 459604 86000
rect 459004 -5282 459186 -5046
rect 459422 -5282 459604 -5046
rect 459004 -5366 459604 -5282
rect 459004 -5602 459186 -5366
rect 459422 -5602 459604 -5366
rect 459004 -5624 459604 -5602
rect 444604 -6222 444786 -5986
rect 445022 -6222 445204 -5986
rect 444604 -6306 445204 -6222
rect 444604 -6542 444786 -6306
rect 445022 -6542 445204 -6306
rect 444604 -7504 445204 -6542
rect 462604 -6926 463204 86000
rect 473404 -2226 474004 86000
rect 473404 -2462 473586 -2226
rect 473822 -2462 474004 -2226
rect 473404 -2546 474004 -2462
rect 473404 -2782 473586 -2546
rect 473822 -2782 474004 -2546
rect 473404 -3744 474004 -2782
rect 477004 -4106 477604 86000
rect 477004 -4342 477186 -4106
rect 477422 -4342 477604 -4106
rect 477004 -4426 477604 -4342
rect 477004 -4662 477186 -4426
rect 477422 -4662 477604 -4426
rect 477004 -5624 477604 -4662
rect 462604 -7162 462786 -6926
rect 463022 -7162 463204 -6926
rect 462604 -7246 463204 -7162
rect 462604 -7482 462786 -7246
rect 463022 -7482 463204 -7246
rect 462604 -7504 463204 -7482
rect 480604 -5986 481204 86000
rect 491404 -3166 492004 86000
rect 491404 -3402 491586 -3166
rect 491822 -3402 492004 -3166
rect 491404 -3486 492004 -3402
rect 491404 -3722 491586 -3486
rect 491822 -3722 492004 -3486
rect 491404 -3744 492004 -3722
rect 495004 -5046 495604 86000
rect 495004 -5282 495186 -5046
rect 495422 -5282 495604 -5046
rect 495004 -5366 495604 -5282
rect 495004 -5602 495186 -5366
rect 495422 -5602 495604 -5366
rect 495004 -5624 495604 -5602
rect 480604 -6222 480786 -5986
rect 481022 -6222 481204 -5986
rect 480604 -6306 481204 -6222
rect 480604 -6542 480786 -6306
rect 481022 -6542 481204 -6306
rect 480604 -7504 481204 -6542
rect 498604 -6926 499204 86000
rect 509404 -2226 510004 86000
rect 509404 -2462 509586 -2226
rect 509822 -2462 510004 -2226
rect 509404 -2546 510004 -2462
rect 509404 -2782 509586 -2546
rect 509822 -2782 510004 -2546
rect 509404 -3744 510004 -2782
rect 513004 -4106 513604 86000
rect 513004 -4342 513186 -4106
rect 513422 -4342 513604 -4106
rect 513004 -4426 513604 -4342
rect 513004 -4662 513186 -4426
rect 513422 -4662 513604 -4426
rect 513004 -5624 513604 -4662
rect 498604 -7162 498786 -6926
rect 499022 -7162 499204 -6926
rect 498604 -7246 499204 -7162
rect 498604 -7482 498786 -7246
rect 499022 -7482 499204 -7246
rect 498604 -7504 499204 -7482
rect 516604 -5986 517204 86000
rect 527404 -3166 528004 707102
rect 527404 -3402 527586 -3166
rect 527822 -3402 528004 -3166
rect 527404 -3486 528004 -3402
rect 527404 -3722 527586 -3486
rect 527822 -3722 528004 -3486
rect 527404 -3744 528004 -3722
rect 531004 -5046 531604 708982
rect 531004 -5282 531186 -5046
rect 531422 -5282 531604 -5046
rect 531004 -5366 531604 -5282
rect 531004 -5602 531186 -5366
rect 531422 -5602 531604 -5366
rect 531004 -5624 531604 -5602
rect 516604 -6222 516786 -5986
rect 517022 -6222 517204 -5986
rect 516604 -6306 517204 -6222
rect 516604 -6542 516786 -6306
rect 517022 -6542 517204 -6306
rect 516604 -7504 517204 -6542
rect 534604 -6926 535204 710862
rect 552604 710478 553204 711440
rect 552604 710242 552786 710478
rect 553022 710242 553204 710478
rect 552604 710158 553204 710242
rect 552604 709922 552786 710158
rect 553022 709922 553204 710158
rect 549004 708598 549604 709560
rect 549004 708362 549186 708598
rect 549422 708362 549604 708598
rect 549004 708278 549604 708362
rect 549004 708042 549186 708278
rect 549422 708042 549604 708278
rect 545404 706718 546004 707680
rect 545404 706482 545586 706718
rect 545822 706482 546004 706718
rect 545404 706398 546004 706482
rect 545404 706162 545586 706398
rect 545822 706162 546004 706398
rect 545404 -2226 546004 706162
rect 545404 -2462 545586 -2226
rect 545822 -2462 546004 -2226
rect 545404 -2546 546004 -2462
rect 545404 -2782 545586 -2546
rect 545822 -2782 546004 -2546
rect 545404 -3744 546004 -2782
rect 549004 -4106 549604 708042
rect 549004 -4342 549186 -4106
rect 549422 -4342 549604 -4106
rect 549004 -4426 549604 -4342
rect 549004 -4662 549186 -4426
rect 549422 -4662 549604 -4426
rect 549004 -5624 549604 -4662
rect 534604 -7162 534786 -6926
rect 535022 -7162 535204 -6926
rect 534604 -7246 535204 -7162
rect 534604 -7482 534786 -7246
rect 535022 -7482 535204 -7246
rect 534604 -7504 535204 -7482
rect 552604 -5986 553204 709922
rect 570604 711418 571204 711440
rect 570604 711182 570786 711418
rect 571022 711182 571204 711418
rect 570604 711098 571204 711182
rect 570604 710862 570786 711098
rect 571022 710862 571204 711098
rect 567004 709538 567604 709560
rect 567004 709302 567186 709538
rect 567422 709302 567604 709538
rect 567004 709218 567604 709302
rect 567004 708982 567186 709218
rect 567422 708982 567604 709218
rect 563404 707658 564004 707680
rect 563404 707422 563586 707658
rect 563822 707422 564004 707658
rect 563404 707338 564004 707422
rect 563404 707102 563586 707338
rect 563822 707102 564004 707338
rect 563404 -3166 564004 707102
rect 563404 -3402 563586 -3166
rect 563822 -3402 564004 -3166
rect 563404 -3486 564004 -3402
rect 563404 -3722 563586 -3486
rect 563822 -3722 564004 -3486
rect 563404 -3744 564004 -3722
rect 567004 -5046 567604 708982
rect 567004 -5282 567186 -5046
rect 567422 -5282 567604 -5046
rect 567004 -5366 567604 -5282
rect 567004 -5602 567186 -5366
rect 567422 -5602 567604 -5366
rect 567004 -5624 567604 -5602
rect 552604 -6222 552786 -5986
rect 553022 -6222 553204 -5986
rect 552604 -6306 553204 -6222
rect 552604 -6542 552786 -6306
rect 553022 -6542 553204 -6306
rect 552604 -7504 553204 -6542
rect 570604 -6926 571204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 581404 706718 582004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 581404 706482 581586 706718
rect 581822 706482 582004 706718
rect 581404 706398 582004 706482
rect 581404 706162 581586 706398
rect 581822 706162 582004 706398
rect 581404 -2226 582004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 692406 585920 704282
rect 585320 692170 585502 692406
rect 585738 692170 585920 692406
rect 585320 692086 585920 692170
rect 585320 691850 585502 692086
rect 585738 691850 585920 692086
rect 585320 677406 585920 691850
rect 585320 677170 585502 677406
rect 585738 677170 585920 677406
rect 585320 677086 585920 677170
rect 585320 676850 585502 677086
rect 585738 676850 585920 677086
rect 585320 662406 585920 676850
rect 585320 662170 585502 662406
rect 585738 662170 585920 662406
rect 585320 662086 585920 662170
rect 585320 661850 585502 662086
rect 585738 661850 585920 662086
rect 585320 -346 585920 661850
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 699906 586860 705222
rect 586260 699670 586442 699906
rect 586678 699670 586860 699906
rect 586260 699586 586860 699670
rect 586260 699350 586442 699586
rect 586678 699350 586860 699586
rect 586260 684906 586860 699350
rect 586260 684670 586442 684906
rect 586678 684670 586860 684906
rect 586260 684586 586860 684670
rect 586260 684350 586442 684586
rect 586678 684350 586860 684586
rect 586260 669906 586860 684350
rect 586260 669670 586442 669906
rect 586678 669670 586860 669906
rect 586260 669586 586860 669670
rect 586260 669350 586442 669586
rect 586678 669350 586860 669586
rect 586260 -1286 586860 669350
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 581404 -2462 581586 -2226
rect 581822 -2462 582004 -2226
rect 581404 -2546 582004 -2462
rect 581404 -2782 581586 -2546
rect 581822 -2782 582004 -2546
rect 581404 -3744 582004 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 570604 -7162 570786 -6926
rect 571022 -7162 571204 -6926
rect 570604 -7246 571204 -7162
rect 570604 -7482 570786 -7246
rect 571022 -7482 571204 -7246
rect 570604 -7504 571204 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 12786 710242 13022 710478
rect 12786 709922 13022 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 9186 708362 9422 708598
rect 9186 708042 9422 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 5586 706482 5822 706718
rect 5586 706162 5822 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 699670 -2518 699906
rect -2754 699350 -2518 699586
rect -2754 684670 -2518 684906
rect -2754 684350 -2518 684586
rect -2754 669670 -2518 669906
rect -2754 669350 -2518 669586
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 692170 -1578 692406
rect -1814 691850 -1578 692086
rect -1814 677170 -1578 677406
rect -1814 676850 -1578 677086
rect -1814 662170 -1578 662406
rect -1814 661850 -1578 662086
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 5586 -2462 5822 -2226
rect 5586 -2782 5822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 9186 -4342 9422 -4106
rect 9186 -4662 9422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 30786 711182 31022 711418
rect 30786 710862 31022 711098
rect 27186 709302 27422 709538
rect 27186 708982 27422 709218
rect 23586 707422 23822 707658
rect 23586 707102 23822 707338
rect 23586 -3402 23822 -3166
rect 23586 -3722 23822 -3486
rect 27186 -5282 27422 -5046
rect 27186 -5602 27422 -5366
rect 12786 -6222 13022 -5986
rect 12786 -6542 13022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 48786 710242 49022 710478
rect 48786 709922 49022 710158
rect 45186 708362 45422 708598
rect 45186 708042 45422 708278
rect 41586 706482 41822 706718
rect 41586 706162 41822 706398
rect 41586 -2462 41822 -2226
rect 41586 -2782 41822 -2546
rect 45186 -4342 45422 -4106
rect 45186 -4662 45422 -4426
rect 30786 -7162 31022 -6926
rect 30786 -7482 31022 -7246
rect 66786 711182 67022 711418
rect 66786 710862 67022 711098
rect 63186 709302 63422 709538
rect 63186 708982 63422 709218
rect 59586 707422 59822 707658
rect 59586 707102 59822 707338
rect 59586 -3402 59822 -3166
rect 59586 -3722 59822 -3486
rect 63186 -5282 63422 -5046
rect 63186 -5602 63422 -5366
rect 48786 -6222 49022 -5986
rect 48786 -6542 49022 -6306
rect 84786 710242 85022 710478
rect 84786 709922 85022 710158
rect 81186 708362 81422 708598
rect 81186 708042 81422 708278
rect 77586 706482 77822 706718
rect 77586 706162 77822 706398
rect 102786 711182 103022 711418
rect 102786 710862 103022 711098
rect 99186 709302 99422 709538
rect 99186 708982 99422 709218
rect 95586 707422 95822 707658
rect 95586 707102 95822 707338
rect 120786 710242 121022 710478
rect 120786 709922 121022 710158
rect 117186 708362 117422 708598
rect 117186 708042 117422 708278
rect 113586 706482 113822 706718
rect 113586 706162 113822 706398
rect 138786 711182 139022 711418
rect 138786 710862 139022 711098
rect 135186 709302 135422 709538
rect 135186 708982 135422 709218
rect 131586 707422 131822 707658
rect 131586 707102 131822 707338
rect 156786 710242 157022 710478
rect 156786 709922 157022 710158
rect 153186 708362 153422 708598
rect 153186 708042 153422 708278
rect 149586 706482 149822 706718
rect 149586 706162 149822 706398
rect 174786 711182 175022 711418
rect 174786 710862 175022 711098
rect 171186 709302 171422 709538
rect 171186 708982 171422 709218
rect 167586 707422 167822 707658
rect 167586 707102 167822 707338
rect 192786 710242 193022 710478
rect 192786 709922 193022 710158
rect 189186 708362 189422 708598
rect 189186 708042 189422 708278
rect 185586 706482 185822 706718
rect 185586 706162 185822 706398
rect 210786 711182 211022 711418
rect 210786 710862 211022 711098
rect 207186 709302 207422 709538
rect 207186 708982 207422 709218
rect 203586 707422 203822 707658
rect 203586 707102 203822 707338
rect 228786 710242 229022 710478
rect 228786 709922 229022 710158
rect 225186 708362 225422 708598
rect 225186 708042 225422 708278
rect 221586 706482 221822 706718
rect 221586 706162 221822 706398
rect 246786 711182 247022 711418
rect 246786 710862 247022 711098
rect 243186 709302 243422 709538
rect 243186 708982 243422 709218
rect 239586 707422 239822 707658
rect 239586 707102 239822 707338
rect 264786 710242 265022 710478
rect 264786 709922 265022 710158
rect 261186 708362 261422 708598
rect 261186 708042 261422 708278
rect 257586 706482 257822 706718
rect 257586 706162 257822 706398
rect 282786 711182 283022 711418
rect 282786 710862 283022 711098
rect 279186 709302 279422 709538
rect 279186 708982 279422 709218
rect 275586 707422 275822 707658
rect 275586 707102 275822 707338
rect 300786 710242 301022 710478
rect 300786 709922 301022 710158
rect 297186 708362 297422 708598
rect 297186 708042 297422 708278
rect 293586 706482 293822 706718
rect 293586 706162 293822 706398
rect 318786 711182 319022 711418
rect 318786 710862 319022 711098
rect 315186 709302 315422 709538
rect 315186 708982 315422 709218
rect 311586 707422 311822 707658
rect 311586 707102 311822 707338
rect 336786 710242 337022 710478
rect 336786 709922 337022 710158
rect 333186 708362 333422 708598
rect 333186 708042 333422 708278
rect 329586 706482 329822 706718
rect 329586 706162 329822 706398
rect 354786 711182 355022 711418
rect 354786 710862 355022 711098
rect 351186 709302 351422 709538
rect 351186 708982 351422 709218
rect 347586 707422 347822 707658
rect 347586 707102 347822 707338
rect 372786 710242 373022 710478
rect 372786 709922 373022 710158
rect 369186 708362 369422 708598
rect 369186 708042 369422 708278
rect 365586 706482 365822 706718
rect 365586 706162 365822 706398
rect 390786 711182 391022 711418
rect 390786 710862 391022 711098
rect 387186 709302 387422 709538
rect 387186 708982 387422 709218
rect 383586 707422 383822 707658
rect 383586 707102 383822 707338
rect 408786 710242 409022 710478
rect 408786 709922 409022 710158
rect 405186 708362 405422 708598
rect 405186 708042 405422 708278
rect 401586 706482 401822 706718
rect 401586 706162 401822 706398
rect 426786 711182 427022 711418
rect 426786 710862 427022 711098
rect 423186 709302 423422 709538
rect 423186 708982 423422 709218
rect 419586 707422 419822 707658
rect 419586 707102 419822 707338
rect 444786 710242 445022 710478
rect 444786 709922 445022 710158
rect 441186 708362 441422 708598
rect 441186 708042 441422 708278
rect 437586 706482 437822 706718
rect 437586 706162 437822 706398
rect 462786 711182 463022 711418
rect 462786 710862 463022 711098
rect 459186 709302 459422 709538
rect 459186 708982 459422 709218
rect 455586 707422 455822 707658
rect 455586 707102 455822 707338
rect 480786 710242 481022 710478
rect 480786 709922 481022 710158
rect 477186 708362 477422 708598
rect 477186 708042 477422 708278
rect 473586 706482 473822 706718
rect 473586 706162 473822 706398
rect 498786 711182 499022 711418
rect 498786 710862 499022 711098
rect 495186 709302 495422 709538
rect 495186 708982 495422 709218
rect 491586 707422 491822 707658
rect 491586 707102 491822 707338
rect 516786 710242 517022 710478
rect 516786 709922 517022 710158
rect 513186 708362 513422 708598
rect 513186 708042 513422 708278
rect 509586 706482 509822 706718
rect 509586 706162 509822 706398
rect 534786 711182 535022 711418
rect 534786 710862 535022 711098
rect 531186 709302 531422 709538
rect 531186 708982 531422 709218
rect 527586 707422 527822 707658
rect 527586 707102 527822 707338
rect 72280 677170 72516 677406
rect 72600 677170 72836 677406
rect 72280 676850 72516 677086
rect 72600 676850 72836 677086
rect 515112 677170 515348 677406
rect 515432 677170 515668 677406
rect 515112 676850 515348 677086
rect 515432 676850 515668 677086
rect 71120 669670 71356 669906
rect 71440 669670 71676 669906
rect 71120 669350 71356 669586
rect 71440 669350 71676 669586
rect 516272 669670 516508 669906
rect 516592 669670 516828 669906
rect 516272 669350 516508 669586
rect 516592 669350 516828 669586
rect 72280 662170 72516 662406
rect 72600 662170 72836 662406
rect 72280 661850 72516 662086
rect 72600 661850 72836 662086
rect 515112 662170 515348 662406
rect 515432 662170 515668 662406
rect 515112 661850 515348 662086
rect 515432 661850 515668 662086
rect 77586 -2462 77822 -2226
rect 77586 -2782 77822 -2546
rect 81186 -4342 81422 -4106
rect 81186 -4662 81422 -4426
rect 66786 -7162 67022 -6926
rect 66786 -7482 67022 -7246
rect 95586 -3402 95822 -3166
rect 95586 -3722 95822 -3486
rect 99186 -5282 99422 -5046
rect 99186 -5602 99422 -5366
rect 84786 -6222 85022 -5986
rect 84786 -6542 85022 -6306
rect 113586 -2462 113822 -2226
rect 113586 -2782 113822 -2546
rect 117186 -4342 117422 -4106
rect 117186 -4662 117422 -4426
rect 102786 -7162 103022 -6926
rect 102786 -7482 103022 -7246
rect 131586 -3402 131822 -3166
rect 131586 -3722 131822 -3486
rect 135186 -5282 135422 -5046
rect 135186 -5602 135422 -5366
rect 120786 -6222 121022 -5986
rect 120786 -6542 121022 -6306
rect 149586 -2462 149822 -2226
rect 149586 -2782 149822 -2546
rect 153186 -4342 153422 -4106
rect 153186 -4662 153422 -4426
rect 138786 -7162 139022 -6926
rect 138786 -7482 139022 -7246
rect 167586 -3402 167822 -3166
rect 167586 -3722 167822 -3486
rect 171186 -5282 171422 -5046
rect 171186 -5602 171422 -5366
rect 156786 -6222 157022 -5986
rect 156786 -6542 157022 -6306
rect 185586 -2462 185822 -2226
rect 185586 -2782 185822 -2546
rect 189186 -4342 189422 -4106
rect 189186 -4662 189422 -4426
rect 174786 -7162 175022 -6926
rect 174786 -7482 175022 -7246
rect 203586 -3402 203822 -3166
rect 203586 -3722 203822 -3486
rect 207186 -5282 207422 -5046
rect 207186 -5602 207422 -5366
rect 192786 -6222 193022 -5986
rect 192786 -6542 193022 -6306
rect 221586 -2462 221822 -2226
rect 221586 -2782 221822 -2546
rect 225186 -4342 225422 -4106
rect 225186 -4662 225422 -4426
rect 210786 -7162 211022 -6926
rect 210786 -7482 211022 -7246
rect 239586 -3402 239822 -3166
rect 239586 -3722 239822 -3486
rect 243186 -5282 243422 -5046
rect 243186 -5602 243422 -5366
rect 228786 -6222 229022 -5986
rect 228786 -6542 229022 -6306
rect 257586 -2462 257822 -2226
rect 257586 -2782 257822 -2546
rect 261186 -4342 261422 -4106
rect 261186 -4662 261422 -4426
rect 246786 -7162 247022 -6926
rect 246786 -7482 247022 -7246
rect 275586 -3402 275822 -3166
rect 275586 -3722 275822 -3486
rect 279186 -5282 279422 -5046
rect 279186 -5602 279422 -5366
rect 264786 -6222 265022 -5986
rect 264786 -6542 265022 -6306
rect 293586 -2462 293822 -2226
rect 293586 -2782 293822 -2546
rect 297186 -4342 297422 -4106
rect 297186 -4662 297422 -4426
rect 282786 -7162 283022 -6926
rect 282786 -7482 283022 -7246
rect 311586 -3402 311822 -3166
rect 311586 -3722 311822 -3486
rect 315186 -5282 315422 -5046
rect 315186 -5602 315422 -5366
rect 300786 -6222 301022 -5986
rect 300786 -6542 301022 -6306
rect 329586 -2462 329822 -2226
rect 329586 -2782 329822 -2546
rect 333186 -4342 333422 -4106
rect 333186 -4662 333422 -4426
rect 318786 -7162 319022 -6926
rect 318786 -7482 319022 -7246
rect 347586 -3402 347822 -3166
rect 347586 -3722 347822 -3486
rect 351186 -5282 351422 -5046
rect 351186 -5602 351422 -5366
rect 336786 -6222 337022 -5986
rect 336786 -6542 337022 -6306
rect 365586 -2462 365822 -2226
rect 365586 -2782 365822 -2546
rect 369186 -4342 369422 -4106
rect 369186 -4662 369422 -4426
rect 354786 -7162 355022 -6926
rect 354786 -7482 355022 -7246
rect 383586 -3402 383822 -3166
rect 383586 -3722 383822 -3486
rect 387186 -5282 387422 -5046
rect 387186 -5602 387422 -5366
rect 372786 -6222 373022 -5986
rect 372786 -6542 373022 -6306
rect 401586 -2462 401822 -2226
rect 401586 -2782 401822 -2546
rect 405186 -4342 405422 -4106
rect 405186 -4662 405422 -4426
rect 390786 -7162 391022 -6926
rect 390786 -7482 391022 -7246
rect 419586 -3402 419822 -3166
rect 419586 -3722 419822 -3486
rect 423186 -5282 423422 -5046
rect 423186 -5602 423422 -5366
rect 408786 -6222 409022 -5986
rect 408786 -6542 409022 -6306
rect 437586 -2462 437822 -2226
rect 437586 -2782 437822 -2546
rect 441186 -4342 441422 -4106
rect 441186 -4662 441422 -4426
rect 426786 -7162 427022 -6926
rect 426786 -7482 427022 -7246
rect 455586 -3402 455822 -3166
rect 455586 -3722 455822 -3486
rect 459186 -5282 459422 -5046
rect 459186 -5602 459422 -5366
rect 444786 -6222 445022 -5986
rect 444786 -6542 445022 -6306
rect 473586 -2462 473822 -2226
rect 473586 -2782 473822 -2546
rect 477186 -4342 477422 -4106
rect 477186 -4662 477422 -4426
rect 462786 -7162 463022 -6926
rect 462786 -7482 463022 -7246
rect 491586 -3402 491822 -3166
rect 491586 -3722 491822 -3486
rect 495186 -5282 495422 -5046
rect 495186 -5602 495422 -5366
rect 480786 -6222 481022 -5986
rect 480786 -6542 481022 -6306
rect 509586 -2462 509822 -2226
rect 509586 -2782 509822 -2546
rect 513186 -4342 513422 -4106
rect 513186 -4662 513422 -4426
rect 498786 -7162 499022 -6926
rect 498786 -7482 499022 -7246
rect 527586 -3402 527822 -3166
rect 527586 -3722 527822 -3486
rect 531186 -5282 531422 -5046
rect 531186 -5602 531422 -5366
rect 516786 -6222 517022 -5986
rect 516786 -6542 517022 -6306
rect 552786 710242 553022 710478
rect 552786 709922 553022 710158
rect 549186 708362 549422 708598
rect 549186 708042 549422 708278
rect 545586 706482 545822 706718
rect 545586 706162 545822 706398
rect 545586 -2462 545822 -2226
rect 545586 -2782 545822 -2546
rect 549186 -4342 549422 -4106
rect 549186 -4662 549422 -4426
rect 534786 -7162 535022 -6926
rect 534786 -7482 535022 -7246
rect 570786 711182 571022 711418
rect 570786 710862 571022 711098
rect 567186 709302 567422 709538
rect 567186 708982 567422 709218
rect 563586 707422 563822 707658
rect 563586 707102 563822 707338
rect 563586 -3402 563822 -3166
rect 563586 -3722 563822 -3486
rect 567186 -5282 567422 -5046
rect 567186 -5602 567422 -5366
rect 552786 -6222 553022 -5986
rect 552786 -6542 553022 -6306
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 581586 706482 581822 706718
rect 581586 706162 581822 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 692170 585738 692406
rect 585502 691850 585738 692086
rect 585502 677170 585738 677406
rect 585502 676850 585738 677086
rect 585502 662170 585738 662406
rect 585502 661850 585738 662086
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 699670 586678 699906
rect 586442 699350 586678 699586
rect 586442 684670 586678 684906
rect 586442 684350 586678 684586
rect 586442 669670 586678 669906
rect 586442 669350 586678 669586
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 581586 -2462 581822 -2226
rect 581586 -2782 581822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 570786 -7162 571022 -6926
rect 570786 -7482 571022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 30786 711418
rect 31022 711182 66786 711418
rect 67022 711182 102786 711418
rect 103022 711182 138786 711418
rect 139022 711182 174786 711418
rect 175022 711182 210786 711418
rect 211022 711182 246786 711418
rect 247022 711182 282786 711418
rect 283022 711182 318786 711418
rect 319022 711182 354786 711418
rect 355022 711182 390786 711418
rect 391022 711182 426786 711418
rect 427022 711182 462786 711418
rect 463022 711182 498786 711418
rect 499022 711182 534786 711418
rect 535022 711182 570786 711418
rect 571022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 30786 711098
rect 31022 710862 66786 711098
rect 67022 710862 102786 711098
rect 103022 710862 138786 711098
rect 139022 710862 174786 711098
rect 175022 710862 210786 711098
rect 211022 710862 246786 711098
rect 247022 710862 282786 711098
rect 283022 710862 318786 711098
rect 319022 710862 354786 711098
rect 355022 710862 390786 711098
rect 391022 710862 426786 711098
rect 427022 710862 462786 711098
rect 463022 710862 498786 711098
rect 499022 710862 534786 711098
rect 535022 710862 570786 711098
rect 571022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 12786 710478
rect 13022 710242 48786 710478
rect 49022 710242 84786 710478
rect 85022 710242 120786 710478
rect 121022 710242 156786 710478
rect 157022 710242 192786 710478
rect 193022 710242 228786 710478
rect 229022 710242 264786 710478
rect 265022 710242 300786 710478
rect 301022 710242 336786 710478
rect 337022 710242 372786 710478
rect 373022 710242 408786 710478
rect 409022 710242 444786 710478
rect 445022 710242 480786 710478
rect 481022 710242 516786 710478
rect 517022 710242 552786 710478
rect 553022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 12786 710158
rect 13022 709922 48786 710158
rect 49022 709922 84786 710158
rect 85022 709922 120786 710158
rect 121022 709922 156786 710158
rect 157022 709922 192786 710158
rect 193022 709922 228786 710158
rect 229022 709922 264786 710158
rect 265022 709922 300786 710158
rect 301022 709922 336786 710158
rect 337022 709922 372786 710158
rect 373022 709922 408786 710158
rect 409022 709922 444786 710158
rect 445022 709922 480786 710158
rect 481022 709922 516786 710158
rect 517022 709922 552786 710158
rect 553022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 27186 709538
rect 27422 709302 63186 709538
rect 63422 709302 99186 709538
rect 99422 709302 135186 709538
rect 135422 709302 171186 709538
rect 171422 709302 207186 709538
rect 207422 709302 243186 709538
rect 243422 709302 279186 709538
rect 279422 709302 315186 709538
rect 315422 709302 351186 709538
rect 351422 709302 387186 709538
rect 387422 709302 423186 709538
rect 423422 709302 459186 709538
rect 459422 709302 495186 709538
rect 495422 709302 531186 709538
rect 531422 709302 567186 709538
rect 567422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 27186 709218
rect 27422 708982 63186 709218
rect 63422 708982 99186 709218
rect 99422 708982 135186 709218
rect 135422 708982 171186 709218
rect 171422 708982 207186 709218
rect 207422 708982 243186 709218
rect 243422 708982 279186 709218
rect 279422 708982 315186 709218
rect 315422 708982 351186 709218
rect 351422 708982 387186 709218
rect 387422 708982 423186 709218
rect 423422 708982 459186 709218
rect 459422 708982 495186 709218
rect 495422 708982 531186 709218
rect 531422 708982 567186 709218
rect 567422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 9186 708598
rect 9422 708362 45186 708598
rect 45422 708362 81186 708598
rect 81422 708362 117186 708598
rect 117422 708362 153186 708598
rect 153422 708362 189186 708598
rect 189422 708362 225186 708598
rect 225422 708362 261186 708598
rect 261422 708362 297186 708598
rect 297422 708362 333186 708598
rect 333422 708362 369186 708598
rect 369422 708362 405186 708598
rect 405422 708362 441186 708598
rect 441422 708362 477186 708598
rect 477422 708362 513186 708598
rect 513422 708362 549186 708598
rect 549422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 9186 708278
rect 9422 708042 45186 708278
rect 45422 708042 81186 708278
rect 81422 708042 117186 708278
rect 117422 708042 153186 708278
rect 153422 708042 189186 708278
rect 189422 708042 225186 708278
rect 225422 708042 261186 708278
rect 261422 708042 297186 708278
rect 297422 708042 333186 708278
rect 333422 708042 369186 708278
rect 369422 708042 405186 708278
rect 405422 708042 441186 708278
rect 441422 708042 477186 708278
rect 477422 708042 513186 708278
rect 513422 708042 549186 708278
rect 549422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 23586 707658
rect 23822 707422 59586 707658
rect 59822 707422 95586 707658
rect 95822 707422 131586 707658
rect 131822 707422 167586 707658
rect 167822 707422 203586 707658
rect 203822 707422 239586 707658
rect 239822 707422 275586 707658
rect 275822 707422 311586 707658
rect 311822 707422 347586 707658
rect 347822 707422 383586 707658
rect 383822 707422 419586 707658
rect 419822 707422 455586 707658
rect 455822 707422 491586 707658
rect 491822 707422 527586 707658
rect 527822 707422 563586 707658
rect 563822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 23586 707338
rect 23822 707102 59586 707338
rect 59822 707102 95586 707338
rect 95822 707102 131586 707338
rect 131822 707102 167586 707338
rect 167822 707102 203586 707338
rect 203822 707102 239586 707338
rect 239822 707102 275586 707338
rect 275822 707102 311586 707338
rect 311822 707102 347586 707338
rect 347822 707102 383586 707338
rect 383822 707102 419586 707338
rect 419822 707102 455586 707338
rect 455822 707102 491586 707338
rect 491822 707102 527586 707338
rect 527822 707102 563586 707338
rect 563822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 5586 706718
rect 5822 706482 41586 706718
rect 41822 706482 77586 706718
rect 77822 706482 113586 706718
rect 113822 706482 149586 706718
rect 149822 706482 185586 706718
rect 185822 706482 221586 706718
rect 221822 706482 257586 706718
rect 257822 706482 293586 706718
rect 293822 706482 329586 706718
rect 329822 706482 365586 706718
rect 365822 706482 401586 706718
rect 401822 706482 437586 706718
rect 437822 706482 473586 706718
rect 473822 706482 509586 706718
rect 509822 706482 545586 706718
rect 545822 706482 581586 706718
rect 581822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 5586 706398
rect 5822 706162 41586 706398
rect 41822 706162 77586 706398
rect 77822 706162 113586 706398
rect 113822 706162 149586 706398
rect 149822 706162 185586 706398
rect 185822 706162 221586 706398
rect 221822 706162 257586 706398
rect 257822 706162 293586 706398
rect 293822 706162 329586 706398
rect 329822 706162 365586 706398
rect 365822 706162 401586 706398
rect 401822 706162 437586 706398
rect 437822 706162 473586 706398
rect 473822 706162 509586 706398
rect 509822 706162 545586 706398
rect 545822 706162 581586 706398
rect 581822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 585320 704258 585920 704260
rect -2936 699928 -2336 699930
rect 586260 699928 586860 699930
rect -2936 699906 586860 699928
rect -2936 699670 -2754 699906
rect -2518 699670 586442 699906
rect 586678 699670 586860 699906
rect -2936 699586 586860 699670
rect -2936 699350 -2754 699586
rect -2518 699350 586442 699586
rect 586678 699350 586860 699586
rect -2936 699328 586860 699350
rect -2936 699326 -2336 699328
rect 586260 699326 586860 699328
rect -1996 692428 -1396 692430
rect 585320 692428 585920 692430
rect -2936 692406 586860 692428
rect -2936 692170 -1814 692406
rect -1578 692170 585502 692406
rect 585738 692170 586860 692406
rect -2936 692086 586860 692170
rect -2936 691850 -1814 692086
rect -1578 691850 585502 692086
rect 585738 691850 586860 692086
rect -2936 691828 586860 691850
rect -1996 691826 -1396 691828
rect 585320 691826 585920 691828
rect -2936 684928 -2336 684930
rect 586260 684928 586860 684930
rect -2936 684906 586860 684928
rect -2936 684670 -2754 684906
rect -2518 684670 586442 684906
rect 586678 684670 586860 684906
rect -2936 684586 586860 684670
rect -2936 684350 -2754 684586
rect -2518 684350 586442 684586
rect 586678 684350 586860 684586
rect -2936 684328 586860 684350
rect -2936 684326 -2336 684328
rect 586260 684326 586860 684328
rect -1996 677428 -1396 677430
rect 72158 677428 72958 677430
rect 514990 677428 515790 677430
rect 585320 677428 585920 677430
rect -2936 677406 586860 677428
rect -2936 677170 -1814 677406
rect -1578 677170 72280 677406
rect 72516 677170 72600 677406
rect 72836 677170 515112 677406
rect 515348 677170 515432 677406
rect 515668 677170 585502 677406
rect 585738 677170 586860 677406
rect -2936 677086 586860 677170
rect -2936 676850 -1814 677086
rect -1578 676850 72280 677086
rect 72516 676850 72600 677086
rect 72836 676850 515112 677086
rect 515348 676850 515432 677086
rect 515668 676850 585502 677086
rect 585738 676850 586860 677086
rect -2936 676828 586860 676850
rect -1996 676826 -1396 676828
rect 72158 676826 72958 676828
rect 514990 676826 515790 676828
rect 585320 676826 585920 676828
rect -2936 669928 -2336 669930
rect 70998 669928 71798 669930
rect 516150 669928 516950 669930
rect 586260 669928 586860 669930
rect -2936 669906 586860 669928
rect -2936 669670 -2754 669906
rect -2518 669670 71120 669906
rect 71356 669670 71440 669906
rect 71676 669670 516272 669906
rect 516508 669670 516592 669906
rect 516828 669670 586442 669906
rect 586678 669670 586860 669906
rect -2936 669586 586860 669670
rect -2936 669350 -2754 669586
rect -2518 669350 71120 669586
rect 71356 669350 71440 669586
rect 71676 669350 516272 669586
rect 516508 669350 516592 669586
rect 516828 669350 586442 669586
rect 586678 669350 586860 669586
rect -2936 669328 586860 669350
rect -2936 669326 -2336 669328
rect 70998 669326 71798 669328
rect 516150 669326 516950 669328
rect 586260 669326 586860 669328
rect -1996 662428 -1396 662430
rect 72158 662428 72958 662430
rect 514990 662428 515790 662430
rect 585320 662428 585920 662430
rect -2936 662406 586860 662428
rect -2936 662170 -1814 662406
rect -1578 662170 72280 662406
rect 72516 662170 72600 662406
rect 72836 662170 515112 662406
rect 515348 662170 515432 662406
rect 515668 662170 585502 662406
rect 585738 662170 586860 662406
rect -2936 662086 586860 662170
rect -2936 661850 -1814 662086
rect -1578 661850 72280 662086
rect 72516 661850 72600 662086
rect 72836 661850 515112 662086
rect 515348 661850 515432 662086
rect 515668 661850 585502 662086
rect 585738 661850 586860 662086
rect -2936 661828 586860 661850
rect -1996 661826 -1396 661828
rect 72158 661826 72958 661828
rect 514990 661826 515790 661828
rect 585320 661826 585920 661828
rect -1996 -324 -1396 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 5586 -2226
rect 5822 -2462 41586 -2226
rect 41822 -2462 77586 -2226
rect 77822 -2462 113586 -2226
rect 113822 -2462 149586 -2226
rect 149822 -2462 185586 -2226
rect 185822 -2462 221586 -2226
rect 221822 -2462 257586 -2226
rect 257822 -2462 293586 -2226
rect 293822 -2462 329586 -2226
rect 329822 -2462 365586 -2226
rect 365822 -2462 401586 -2226
rect 401822 -2462 437586 -2226
rect 437822 -2462 473586 -2226
rect 473822 -2462 509586 -2226
rect 509822 -2462 545586 -2226
rect 545822 -2462 581586 -2226
rect 581822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 5586 -2546
rect 5822 -2782 41586 -2546
rect 41822 -2782 77586 -2546
rect 77822 -2782 113586 -2546
rect 113822 -2782 149586 -2546
rect 149822 -2782 185586 -2546
rect 185822 -2782 221586 -2546
rect 221822 -2782 257586 -2546
rect 257822 -2782 293586 -2546
rect 293822 -2782 329586 -2546
rect 329822 -2782 365586 -2546
rect 365822 -2782 401586 -2546
rect 401822 -2782 437586 -2546
rect 437822 -2782 473586 -2546
rect 473822 -2782 509586 -2546
rect 509822 -2782 545586 -2546
rect 545822 -2782 581586 -2546
rect 581822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 23586 -3166
rect 23822 -3402 59586 -3166
rect 59822 -3402 95586 -3166
rect 95822 -3402 131586 -3166
rect 131822 -3402 167586 -3166
rect 167822 -3402 203586 -3166
rect 203822 -3402 239586 -3166
rect 239822 -3402 275586 -3166
rect 275822 -3402 311586 -3166
rect 311822 -3402 347586 -3166
rect 347822 -3402 383586 -3166
rect 383822 -3402 419586 -3166
rect 419822 -3402 455586 -3166
rect 455822 -3402 491586 -3166
rect 491822 -3402 527586 -3166
rect 527822 -3402 563586 -3166
rect 563822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 23586 -3486
rect 23822 -3722 59586 -3486
rect 59822 -3722 95586 -3486
rect 95822 -3722 131586 -3486
rect 131822 -3722 167586 -3486
rect 167822 -3722 203586 -3486
rect 203822 -3722 239586 -3486
rect 239822 -3722 275586 -3486
rect 275822 -3722 311586 -3486
rect 311822 -3722 347586 -3486
rect 347822 -3722 383586 -3486
rect 383822 -3722 419586 -3486
rect 419822 -3722 455586 -3486
rect 455822 -3722 491586 -3486
rect 491822 -3722 527586 -3486
rect 527822 -3722 563586 -3486
rect 563822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 9186 -4106
rect 9422 -4342 45186 -4106
rect 45422 -4342 81186 -4106
rect 81422 -4342 117186 -4106
rect 117422 -4342 153186 -4106
rect 153422 -4342 189186 -4106
rect 189422 -4342 225186 -4106
rect 225422 -4342 261186 -4106
rect 261422 -4342 297186 -4106
rect 297422 -4342 333186 -4106
rect 333422 -4342 369186 -4106
rect 369422 -4342 405186 -4106
rect 405422 -4342 441186 -4106
rect 441422 -4342 477186 -4106
rect 477422 -4342 513186 -4106
rect 513422 -4342 549186 -4106
rect 549422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 9186 -4426
rect 9422 -4662 45186 -4426
rect 45422 -4662 81186 -4426
rect 81422 -4662 117186 -4426
rect 117422 -4662 153186 -4426
rect 153422 -4662 189186 -4426
rect 189422 -4662 225186 -4426
rect 225422 -4662 261186 -4426
rect 261422 -4662 297186 -4426
rect 297422 -4662 333186 -4426
rect 333422 -4662 369186 -4426
rect 369422 -4662 405186 -4426
rect 405422 -4662 441186 -4426
rect 441422 -4662 477186 -4426
rect 477422 -4662 513186 -4426
rect 513422 -4662 549186 -4426
rect 549422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 27186 -5046
rect 27422 -5282 63186 -5046
rect 63422 -5282 99186 -5046
rect 99422 -5282 135186 -5046
rect 135422 -5282 171186 -5046
rect 171422 -5282 207186 -5046
rect 207422 -5282 243186 -5046
rect 243422 -5282 279186 -5046
rect 279422 -5282 315186 -5046
rect 315422 -5282 351186 -5046
rect 351422 -5282 387186 -5046
rect 387422 -5282 423186 -5046
rect 423422 -5282 459186 -5046
rect 459422 -5282 495186 -5046
rect 495422 -5282 531186 -5046
rect 531422 -5282 567186 -5046
rect 567422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 27186 -5366
rect 27422 -5602 63186 -5366
rect 63422 -5602 99186 -5366
rect 99422 -5602 135186 -5366
rect 135422 -5602 171186 -5366
rect 171422 -5602 207186 -5366
rect 207422 -5602 243186 -5366
rect 243422 -5602 279186 -5366
rect 279422 -5602 315186 -5366
rect 315422 -5602 351186 -5366
rect 351422 -5602 387186 -5366
rect 387422 -5602 423186 -5366
rect 423422 -5602 459186 -5366
rect 459422 -5602 495186 -5366
rect 495422 -5602 531186 -5366
rect 531422 -5602 567186 -5366
rect 567422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 12786 -5986
rect 13022 -6222 48786 -5986
rect 49022 -6222 84786 -5986
rect 85022 -6222 120786 -5986
rect 121022 -6222 156786 -5986
rect 157022 -6222 192786 -5986
rect 193022 -6222 228786 -5986
rect 229022 -6222 264786 -5986
rect 265022 -6222 300786 -5986
rect 301022 -6222 336786 -5986
rect 337022 -6222 372786 -5986
rect 373022 -6222 408786 -5986
rect 409022 -6222 444786 -5986
rect 445022 -6222 480786 -5986
rect 481022 -6222 516786 -5986
rect 517022 -6222 552786 -5986
rect 553022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 12786 -6306
rect 13022 -6542 48786 -6306
rect 49022 -6542 84786 -6306
rect 85022 -6542 120786 -6306
rect 121022 -6542 156786 -6306
rect 157022 -6542 192786 -6306
rect 193022 -6542 228786 -6306
rect 229022 -6542 264786 -6306
rect 265022 -6542 300786 -6306
rect 301022 -6542 336786 -6306
rect 337022 -6542 372786 -6306
rect 373022 -6542 408786 -6306
rect 409022 -6542 444786 -6306
rect 445022 -6542 480786 -6306
rect 481022 -6542 516786 -6306
rect 517022 -6542 552786 -6306
rect 553022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 30786 -6926
rect 31022 -7162 66786 -6926
rect 67022 -7162 102786 -6926
rect 103022 -7162 138786 -6926
rect 139022 -7162 174786 -6926
rect 175022 -7162 210786 -6926
rect 211022 -7162 246786 -6926
rect 247022 -7162 282786 -6926
rect 283022 -7162 318786 -6926
rect 319022 -7162 354786 -6926
rect 355022 -7162 390786 -6926
rect 391022 -7162 426786 -6926
rect 427022 -7162 462786 -6926
rect 463022 -7162 498786 -6926
rect 499022 -7162 534786 -6926
rect 535022 -7162 570786 -6926
rect 571022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 30786 -7246
rect 31022 -7482 66786 -7246
rect 67022 -7482 102786 -7246
rect 103022 -7482 138786 -7246
rect 139022 -7482 174786 -7246
rect 175022 -7482 210786 -7246
rect 211022 -7482 246786 -7246
rect 247022 -7482 282786 -7246
rect 283022 -7482 318786 -7246
rect 319022 -7482 354786 -7246
rect 355022 -7482 390786 -7246
rect 391022 -7482 426786 -7246
rect 427022 -7482 462786 -7246
rect 463022 -7482 498786 -7246
rect 499022 -7482 534786 -7246
rect 535022 -7482 570786 -7246
rect 571022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1625000815
transform 1 0 70000 0 1 88000
box 0 0 447948 592008
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 533 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 599 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 600 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 601 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 602 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 603 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 604 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 605 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 606 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 607 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 608 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 609 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 610 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 611 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 612 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 613 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 614 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 615 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 616 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 617 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 618 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 619 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 620 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 621 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 622 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 623 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 624 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 625 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 626 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 627 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 628 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 629 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 630 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1.extra1
port 638 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1.extra2
port 639 nsew power bidirectional
rlabel metal5 s -2936 691828 586860 692428 6 vccd1.extra3
port 640 nsew power bidirectional
rlabel metal5 s -2936 676828 586860 677428 6 vccd1.extra4
port 641 nsew power bidirectional
rlabel metal5 s -2936 661828 586860 662428 6 vccd1.extra5
port 642 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1.extra6
port 643 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 644 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1.extra1
port 645 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1.extra2
port 646 nsew ground bidirectional
rlabel metal5 s -2936 699328 586860 699928 6 vssd1.extra3
port 647 nsew ground bidirectional
rlabel metal5 s -2936 684328 586860 684928 6 vssd1.extra4
port 648 nsew ground bidirectional
rlabel metal5 s -2936 669328 586860 669928 6 vssd1.extra5
port 649 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1.extra6
port 650 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 651 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 707680 6 vccd2.extra1
port 652 nsew power bidirectional
rlabel metal4 s 509404 682008 510004 707680 6 vccd2.extra2
port 653 nsew power bidirectional
rlabel metal4 s 473404 682008 474004 707680 6 vccd2.extra3
port 654 nsew power bidirectional
rlabel metal4 s 437404 682008 438004 707680 6 vccd2.extra4
port 655 nsew power bidirectional
rlabel metal4 s 401404 682008 402004 707680 6 vccd2.extra5
port 656 nsew power bidirectional
rlabel metal4 s 365404 682008 366004 707680 6 vccd2.extra6
port 657 nsew power bidirectional
rlabel metal4 s 329404 682008 330004 707680 6 vccd2.extra7
port 658 nsew power bidirectional
rlabel metal4 s 293404 682008 294004 707680 6 vccd2.extra8
port 659 nsew power bidirectional
rlabel metal4 s 257404 682008 258004 707680 6 vccd2.extra9
port 660 nsew power bidirectional
rlabel metal4 s 221404 682008 222004 707680 6 vccd2.extra10
port 661 nsew power bidirectional
rlabel metal4 s 185404 682008 186004 707680 6 vccd2.extra11
port 662 nsew power bidirectional
rlabel metal4 s 149404 682008 150004 707680 6 vccd2.extra12
port 663 nsew power bidirectional
rlabel metal4 s 113404 682008 114004 707680 6 vccd2.extra13
port 664 nsew power bidirectional
rlabel metal4 s 77404 682008 78004 707680 6 vccd2.extra14
port 665 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 707680 6 vccd2.extra15
port 666 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2.extra16
port 667 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2.extra17
port 668 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2.extra18
port 669 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 86000 6 vccd2.extra19
port 670 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 86000 6 vccd2.extra20
port 671 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 86000 6 vccd2.extra21
port 672 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 86000 6 vccd2.extra22
port 673 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 86000 6 vccd2.extra23
port 674 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 86000 6 vccd2.extra24
port 675 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 86000 6 vccd2.extra25
port 676 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 86000 6 vccd2.extra26
port 677 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 86000 6 vccd2.extra27
port 678 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 86000 6 vccd2.extra28
port 679 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 86000 6 vccd2.extra29
port 680 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 86000 6 vccd2.extra30
port 681 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 86000 6 vccd2.extra31
port 682 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2.extra32
port 683 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2.extra33
port 684 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 685 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 707680 6 vssd2.extra1
port 686 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 707680 6 vssd2.extra2
port 687 nsew ground bidirectional
rlabel metal4 s 491404 682008 492004 707680 6 vssd2.extra3
port 688 nsew ground bidirectional
rlabel metal4 s 455404 682008 456004 707680 6 vssd2.extra4
port 689 nsew ground bidirectional
rlabel metal4 s 419404 682008 420004 707680 6 vssd2.extra5
port 690 nsew ground bidirectional
rlabel metal4 s 383404 682008 384004 707680 6 vssd2.extra6
port 691 nsew ground bidirectional
rlabel metal4 s 347404 682008 348004 707680 6 vssd2.extra7
port 692 nsew ground bidirectional
rlabel metal4 s 311404 682008 312004 707680 6 vssd2.extra8
port 693 nsew ground bidirectional
rlabel metal4 s 275404 682008 276004 707680 6 vssd2.extra9
port 694 nsew ground bidirectional
rlabel metal4 s 239404 682008 240004 707680 6 vssd2.extra10
port 695 nsew ground bidirectional
rlabel metal4 s 203404 682008 204004 707680 6 vssd2.extra11
port 696 nsew ground bidirectional
rlabel metal4 s 167404 682008 168004 707680 6 vssd2.extra12
port 697 nsew ground bidirectional
rlabel metal4 s 131404 682008 132004 707680 6 vssd2.extra13
port 698 nsew ground bidirectional
rlabel metal4 s 95404 682008 96004 707680 6 vssd2.extra14
port 699 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 707680 6 vssd2.extra15
port 700 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2.extra16
port 701 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2.extra17
port 702 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 86000 6 vssd2.extra18
port 703 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 86000 6 vssd2.extra19
port 704 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 86000 6 vssd2.extra20
port 705 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 86000 6 vssd2.extra21
port 706 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 86000 6 vssd2.extra22
port 707 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 86000 6 vssd2.extra23
port 708 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 86000 6 vssd2.extra24
port 709 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 86000 6 vssd2.extra25
port 710 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 86000 6 vssd2.extra26
port 711 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 86000 6 vssd2.extra27
port 712 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 86000 6 vssd2.extra28
port 713 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 86000 6 vssd2.extra29
port 714 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2.extra30
port 715 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2.extra31
port 716 nsew ground bidirectional
rlabel metal4 s 549004 -5624 549604 709560 6 vdda1
port 717 nsew power bidirectional
rlabel metal4 s 513004 682008 513604 709560 6 vdda1.extra1
port 718 nsew power bidirectional
rlabel metal4 s 477004 682008 477604 709560 6 vdda1.extra2
port 719 nsew power bidirectional
rlabel metal4 s 441004 682008 441604 709560 6 vdda1.extra3
port 720 nsew power bidirectional
rlabel metal4 s 405004 682008 405604 709560 6 vdda1.extra4
port 721 nsew power bidirectional
rlabel metal4 s 369004 682008 369604 709560 6 vdda1.extra5
port 722 nsew power bidirectional
rlabel metal4 s 333004 682008 333604 709560 6 vdda1.extra6
port 723 nsew power bidirectional
rlabel metal4 s 297004 682008 297604 709560 6 vdda1.extra7
port 724 nsew power bidirectional
rlabel metal4 s 261004 682008 261604 709560 6 vdda1.extra8
port 725 nsew power bidirectional
rlabel metal4 s 225004 682008 225604 709560 6 vdda1.extra9
port 726 nsew power bidirectional
rlabel metal4 s 189004 682008 189604 709560 6 vdda1.extra10
port 727 nsew power bidirectional
rlabel metal4 s 153004 682008 153604 709560 6 vdda1.extra11
port 728 nsew power bidirectional
rlabel metal4 s 117004 682008 117604 709560 6 vdda1.extra12
port 729 nsew power bidirectional
rlabel metal4 s 81004 682008 81604 709560 6 vdda1.extra13
port 730 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 709560 6 vdda1.extra14
port 731 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1.extra15
port 732 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1.extra16
port 733 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1.extra17
port 734 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 86000 6 vdda1.extra18
port 735 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 86000 6 vdda1.extra19
port 736 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 86000 6 vdda1.extra20
port 737 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 86000 6 vdda1.extra21
port 738 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 86000 6 vdda1.extra22
port 739 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 86000 6 vdda1.extra23
port 740 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 86000 6 vdda1.extra24
port 741 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 86000 6 vdda1.extra25
port 742 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 86000 6 vdda1.extra26
port 743 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 86000 6 vdda1.extra27
port 744 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 86000 6 vdda1.extra28
port 745 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 86000 6 vdda1.extra29
port 746 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 86000 6 vdda1.extra30
port 747 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1.extra31
port 748 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1.extra32
port 749 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 750 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1.extra1
port 751 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 709560 6 vssa1.extra2
port 752 nsew ground bidirectional
rlabel metal4 s 495004 682008 495604 709560 6 vssa1.extra3
port 753 nsew ground bidirectional
rlabel metal4 s 459004 682008 459604 709560 6 vssa1.extra4
port 754 nsew ground bidirectional
rlabel metal4 s 423004 682008 423604 709560 6 vssa1.extra5
port 755 nsew ground bidirectional
rlabel metal4 s 387004 682008 387604 709560 6 vssa1.extra6
port 756 nsew ground bidirectional
rlabel metal4 s 351004 682008 351604 709560 6 vssa1.extra7
port 757 nsew ground bidirectional
rlabel metal4 s 315004 682008 315604 709560 6 vssa1.extra8
port 758 nsew ground bidirectional
rlabel metal4 s 279004 682008 279604 709560 6 vssa1.extra9
port 759 nsew ground bidirectional
rlabel metal4 s 243004 682008 243604 709560 6 vssa1.extra10
port 760 nsew ground bidirectional
rlabel metal4 s 207004 682008 207604 709560 6 vssa1.extra11
port 761 nsew ground bidirectional
rlabel metal4 s 171004 682008 171604 709560 6 vssa1.extra12
port 762 nsew ground bidirectional
rlabel metal4 s 135004 682008 135604 709560 6 vssa1.extra13
port 763 nsew ground bidirectional
rlabel metal4 s 99004 682008 99604 709560 6 vssa1.extra14
port 764 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 709560 6 vssa1.extra15
port 765 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1.extra16
port 766 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1.extra17
port 767 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 86000 6 vssa1.extra18
port 768 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 86000 6 vssa1.extra19
port 769 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 86000 6 vssa1.extra20
port 770 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 86000 6 vssa1.extra21
port 771 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 86000 6 vssa1.extra22
port 772 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 86000 6 vssa1.extra23
port 773 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 86000 6 vssa1.extra24
port 774 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 86000 6 vssa1.extra25
port 775 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 86000 6 vssa1.extra26
port 776 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 86000 6 vssa1.extra27
port 777 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 86000 6 vssa1.extra28
port 778 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 86000 6 vssa1.extra29
port 779 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1.extra30
port 780 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1.extra31
port 781 nsew ground bidirectional
rlabel metal4 s 552604 -7504 553204 711440 6 vdda2
port 782 nsew power bidirectional
rlabel metal4 s 516604 682008 517204 711440 6 vdda2.extra1
port 783 nsew power bidirectional
rlabel metal4 s 480604 682008 481204 711440 6 vdda2.extra2
port 784 nsew power bidirectional
rlabel metal4 s 444604 682008 445204 711440 6 vdda2.extra3
port 785 nsew power bidirectional
rlabel metal4 s 408604 682008 409204 711440 6 vdda2.extra4
port 786 nsew power bidirectional
rlabel metal4 s 372604 682008 373204 711440 6 vdda2.extra5
port 787 nsew power bidirectional
rlabel metal4 s 336604 682008 337204 711440 6 vdda2.extra6
port 788 nsew power bidirectional
rlabel metal4 s 300604 682008 301204 711440 6 vdda2.extra7
port 789 nsew power bidirectional
rlabel metal4 s 264604 682008 265204 711440 6 vdda2.extra8
port 790 nsew power bidirectional
rlabel metal4 s 228604 682008 229204 711440 6 vdda2.extra9
port 791 nsew power bidirectional
rlabel metal4 s 192604 682008 193204 711440 6 vdda2.extra10
port 792 nsew power bidirectional
rlabel metal4 s 156604 682008 157204 711440 6 vdda2.extra11
port 793 nsew power bidirectional
rlabel metal4 s 120604 682008 121204 711440 6 vdda2.extra12
port 794 nsew power bidirectional
rlabel metal4 s 84604 682008 85204 711440 6 vdda2.extra13
port 795 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 711440 6 vdda2.extra14
port 796 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2.extra15
port 797 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2.extra16
port 798 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2.extra17
port 799 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 86000 6 vdda2.extra18
port 800 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 86000 6 vdda2.extra19
port 801 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 86000 6 vdda2.extra20
port 802 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 86000 6 vdda2.extra21
port 803 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 86000 6 vdda2.extra22
port 804 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 86000 6 vdda2.extra23
port 805 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 86000 6 vdda2.extra24
port 806 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 86000 6 vdda2.extra25
port 807 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 86000 6 vdda2.extra26
port 808 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 86000 6 vdda2.extra27
port 809 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 86000 6 vdda2.extra28
port 810 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 86000 6 vdda2.extra29
port 811 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 86000 6 vdda2.extra30
port 812 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2.extra31
port 813 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2.extra32
port 814 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 815 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2.extra1
port 816 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 711440 6 vssa2.extra2
port 817 nsew ground bidirectional
rlabel metal4 s 498604 682008 499204 711440 6 vssa2.extra3
port 818 nsew ground bidirectional
rlabel metal4 s 462604 682008 463204 711440 6 vssa2.extra4
port 819 nsew ground bidirectional
rlabel metal4 s 426604 682008 427204 711440 6 vssa2.extra5
port 820 nsew ground bidirectional
rlabel metal4 s 390604 682008 391204 711440 6 vssa2.extra6
port 821 nsew ground bidirectional
rlabel metal4 s 354604 682008 355204 711440 6 vssa2.extra7
port 822 nsew ground bidirectional
rlabel metal4 s 318604 682008 319204 711440 6 vssa2.extra8
port 823 nsew ground bidirectional
rlabel metal4 s 282604 682008 283204 711440 6 vssa2.extra9
port 824 nsew ground bidirectional
rlabel metal4 s 246604 682008 247204 711440 6 vssa2.extra10
port 825 nsew ground bidirectional
rlabel metal4 s 210604 682008 211204 711440 6 vssa2.extra11
port 826 nsew ground bidirectional
rlabel metal4 s 174604 682008 175204 711440 6 vssa2.extra12
port 827 nsew ground bidirectional
rlabel metal4 s 138604 682008 139204 711440 6 vssa2.extra13
port 828 nsew ground bidirectional
rlabel metal4 s 102604 682008 103204 711440 6 vssa2.extra14
port 829 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 711440 6 vssa2.extra15
port 830 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2.extra16
port 831 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2.extra17
port 832 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 86000 6 vssa2.extra18
port 833 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 86000 6 vssa2.extra19
port 834 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 86000 6 vssa2.extra20
port 835 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 86000 6 vssa2.extra21
port 836 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 86000 6 vssa2.extra22
port 837 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 86000 6 vssa2.extra23
port 838 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 86000 6 vssa2.extra24
port 839 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 86000 6 vssa2.extra25
port 840 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 86000 6 vssa2.extra26
port 841 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 86000 6 vssa2.extra27
port 842 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 86000 6 vssa2.extra28
port 843 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 86000 6 vssa2.extra29
port 844 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2.extra30
port 845 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2.extra31
port 846 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
